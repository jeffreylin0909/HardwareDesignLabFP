module Top(clk, rst, PS2_DATA, PS2_CLK, vgaRed, vgaBlue, vgaGreen, hsync, vsync);
    
    parameter [8:0] A_CODE  = {1'b0, 8'h1C};
    parameter [8:0] D_CODE  = {1'b0, 8'h23};
    parameter [8:0] W_CODE  = {1'b0, 8'h1D};
    parameter [8:0] S_CODE  = {1'b0, 8'h1B};
    
	input clk, rst;//button
	inout PS2_DATA, PS2_CLK;
    output [3:0] vgaRed, vgaGreen, vgaBlue;
    output hsync, vsync;
	
	wire clk_d2;//25MHz
    wire clk_d22;
    wire [16:0] pixel_addr, pixel_addr_m;
    wire [11:0] pixel, pixel_m, RGB_link, RGB_m;
	wire [11:0] data;
    wire valid;
	//640*480
    wire [9:0] h_cnt, v_cnt;
	wire [9:0] h_cnt_re, v_cnt_re;
	
	wire [9:0] pos_h, pos_v;
	
	wire [9:0] pos_h_m, pos_v_m;
	//signals
	wire rst_db;
	wire rst_op;
	
	assign h_cnt_re = h_cnt>>1;
	assign v_cnt_re = v_cnt>>1;
	
	assign RGB_link = (valid==1'b1 && (h_cnt_re+pos_h)%320 < 20 && (v_cnt_re+pos_v)%240 < 20 ) ? pixel : 12'h0;
	assign RGB_m = (valid==1'b1 && (h_cnt_re+pos_h_m)%320 < 20 && (v_cnt_re+pos_v_m)%240 < 20 ) ? pixel_m : 12'h0;
	assign {vgaRed, vgaGreen, vgaBlue} = RGB_link+RGB_m;
	
	//clock
	clk_div #(2) CD0(.clk(clk), .clk_d(clk_d2));
	clk_div #(19) CD1(.clk(clk), .clk_d(clk_d22));
	
	//keyboard
	wire [511:0] key_down;
    wire [8:0] last_change;
    wire been_ready;
	
	//signals
	debounce DB1(.s(rst), .s_db(rst_db), .clk(clk));
	onepulse OP1(.s(rst_db), .s_op(rst_op), .clk(clk_d22));
	
	//control
	state_control SC0(
		.clk(clk_d22),
		.rst(rst_op),
		.A_signal(key_down[A_CODE]),
		.D_signal(key_down[D_CODE]),
		.W_signal(key_down[W_CODE]),
		.S_signal(key_down[S_CODE]),
		.pos_h(pos_h),
		.pos_v(pos_v),
		.pos_h_m(pos_h_m),
		.pos_v_m(pos_v_m)
	);
	mem_addr_gen MAG(
		.h_cnt(h_cnt_re),
		.v_cnt(v_cnt_re), 
		.pos_h(pos_h),
		.pos_v(pos_v),
		.pixel_addr(pixel_addr)
	);
	
	mem_addr_gen MAG_m(
		.h_cnt(h_cnt_re),
		.v_cnt(v_cnt_re), 
		.pos_h(pos_h_m),
		.pos_v(pos_v_m),
		.pixel_addr(pixel_addr_m)
	);
     
	//display
    blk_mem_gen_0 BMG0(
		.clka(clk_d2),
        .wea(0),
        .addra(pixel_addr),
        .dina(data[11:0]),
        .douta(pixel)
    ); 
    
    blk_mem_gen_1 BMG0_m(
		.clka(clk_d2),
        .wea(0),
        .addra(pixel_addr_m),
        .dina(data[11:0]),
        .douta(pixel_m)
    ); 

    vga_controller VC0(
        .pclk(clk_d2),
        .reset(rst),
        .hsync(hsync),
        .vsync(vsync),
        .valid(valid),
        .h_cnt(h_cnt),
        .v_cnt(v_cnt)
    );
	
	KeyboardDecoder key_de (
        .key_down(key_down),
        .last_change(last_change),
        .key_valid(been_ready),
        .PS2_DATA(PS2_DATA),
        .PS2_CLK(PS2_CLK),
        .rst(rst),
        .clk(clk)
    );
	
endmodule