//to generate non-boss stage music
`define NM1 32'd261 //C_freq
`define NM2 32'd277 //C#_freq
`define NM3 32'd294 //D_freq
`define NM4 32'd311 //D#_freq
`define NM5 32'd330 //E_freq
`define NM6 32'd349 //F_freq
`define NM7 32'd370 //F#_freq
`define NM8 32'd392 //G_freq
`define NM9 32'd415 //G#_freq
`define NM10 32'd440 //A_freq
`define NM11 32'd494 //B_freq
`define NM0 32'd20000 //slience (over freq.)

module MusicZelda (
	input [12:0] ibeatNum,	
	output reg [31:0] tone
);
//each block = 1 beat or quarter note
always @(*) begin
	case (ibeatNum)		// 1/16 beat 
		13'd0 : tone = `NM10;	
		13'd1 : tone = `NM10;
		13'd2 : tone = `NM10;
		13'd3 : tone = `NM10;
		13'd4 : tone = `NM10;	
		13'd5 : tone = `NM10;
		13'd6 : tone = `NM10;
		13'd7 : tone = `NM10;
		13'd8 : tone = `NM10;	
		13'd9 : tone = `NM10;
		13'd10 : tone = `NM10;
		13'd11 : tone = `NM10;
		13'd12 : tone = `NM10;	
		13'd13 : tone = `NM10;
		13'd14 : tone = `NM10;
		13'd15 : tone = `NM10;
		
		13'd16 : tone = `NM10;
		13'd17 : tone = `NM10;
		13'd18 : tone = `NM10;
		13'd19 : tone = `NM10;
		13'd20 : tone = `NM10;
		13'd21 : tone = `NM10;
		13'd22 : tone = `NM10;
		13'd23 : tone = `NM10;
		13'd24 : tone = `NM10;
		13'd25 : tone = `NM10;
		13'd26 : tone = `NM10;
		13'd27 : tone = `NM10;
		13'd28 : tone = `NM10;
		13'd29 : tone = `NM10;
		13'd30 : tone = `NM10;
		13'd31 : tone = `NM10;
		
		13'd32 : tone = `NM0;
		13'd33 : tone = `NM0;
		13'd34 : tone = `NM0;
		13'd35 : tone = `NM0;
		13'd36 : tone = `NM0;
		13'd37 : tone = `NM0;
		13'd38 : tone = `NM0;
		13'd39 : tone = `NM0;
		13'd40 : tone = `NM0;
		13'd41 : tone = `NM0;
		13'd42 : tone = `NM0;
		13'd43 : tone = `NM0;
		13'd44 : tone = `NM10;
		13'd45 : tone = `NM10;
		13'd46 : tone = `NM10;
		13'd47 : tone = `NM10;
		
		13'd48 : tone = `NM0;
		13'd49 : tone = `NM10;
		13'd50 : tone = `NM10;
		13'd51 : tone = `NM10;
		13'd52 : tone = `NM10;
		13'd53 : tone = `NM0;
		13'd54 : tone = `NM10;
		13'd55 : tone = `NM10;
		13'd56 : tone = `NM10;
		13'd57 : tone = `NM10;
		13'd58 : tone = `NM0;
		13'd59 : tone = `NM10;
		13'd60 : tone = `NM10;
		13'd61 : tone = `NM10;
		13'd62 : tone = `NM10;
		13'd63 : tone = `NM0;
		
		13'd64 : tone = `NM10;
		13'd65 : tone = `NM10;
		13'd66 : tone = `NM10;
		13'd67 : tone = `NM10;
		13'd68 : tone = `NM10;
		13'd69 : tone = `NM10;
		13'd70 : tone = `NM10;
		13'd71 : tone = `NM10;
		13'd72 : tone = `NM10;
		13'd73 : tone = `NM10;
		13'd74 : tone = `NM10;
		13'd75 : tone = `NM0;
		13'd76 : tone = `NM8;
		13'd77 : tone = `NM8;
		13'd78 : tone = `NM8;
		13'd79 : tone = `NM8;
		
		13'd80 : tone = `NM10;
		13'd81 : tone = `NM10;
		13'd82 : tone = `NM10;
		13'd83 : tone = `NM10;
		13'd84 : tone = `NM10;
		13'd85 : tone = `NM10;
		13'd86 : tone = `NM10;
		13'd87 : tone = `NM10;
		13'd88 : tone = `NM10;
		13'd89 : tone = `NM10;
		13'd90 : tone = `NM10;
		13'd91 : tone = `NM10;
		13'd92 : tone = `NM10;
		13'd93 : tone = `NM10;
		13'd94 : tone = `NM10;
		13'd95 : tone = `NM10;
		
		13'd96 : tone = `NM0;
		13'd97 : tone = `NM0;
		13'd98 : tone = `NM0;
		13'd99 : tone = `NM0;
		13'd100 : tone = `NM0;
		13'd101 : tone = `NM0;
		13'd102 : tone = `NM0;
		13'd103 : tone = `NM0;
		13'd104 : tone = `NM0;
		13'd105 : tone = `NM0;
		13'd106 : tone = `NM0;
		13'd107 : tone = `NM0;
		13'd108 : tone = `NM10;
		13'd109 : tone = `NM10;
		13'd110 : tone = `NM10;
		13'd111 : tone = `NM10;
		
		13'd112 : tone = `NM0;
		13'd113 : tone = `NM10;
		13'd114 : tone = `NM10;
		13'd115 : tone = `NM10;
		13'd116 : tone = `NM10;
		13'd117 : tone = `NM0;
		13'd118 : tone = `NM10;
		13'd119 : tone = `NM10;
		13'd120 : tone = `NM10;
		13'd121 : tone = `NM10;
		13'd122 : tone = `NM0;
		13'd123 : tone = `NM10;
		13'd124 : tone = `NM10;
		13'd125 : tone = `NM10;
		13'd126 : tone = `NM10;
		13'd127 : tone = `NM0;
		
		13'd128 : tone = `NM10;	//3
		13'd129 : tone = `NM10;
		13'd130 : tone = `NM10;
		13'd131 : tone = `NM10;
		13'd132 : tone = `NM10;	//1
		13'd133 : tone = `NM10;
		13'd134 : tone = `NM10;
		13'd135 : tone = `NM10;
		13'd136 : tone = `NM10;	//2
		13'd137 : tone = `NM10;
		13'd138 : tone = `NM10;
		13'd139 : tone = `NM0;
		13'd140 : tone = `NM8;	//6
		13'd141 : tone = `NM8;
		13'd142 : tone = `NM8;
		13'd143 : tone = `NM8;
		
		13'd144 : tone = `NM10;
		13'd145 : tone = `NM10;
		13'd146 : tone = `NM10;
		13'd147 : tone = `NM10;
		13'd148 : tone = `NM10;
		13'd149 : tone = `NM10;
		13'd150 : tone = `NM10;
		13'd151 : tone = `NM10;
		13'd152 : tone = `NM10;
		13'd153 : tone = `NM10;
		13'd154 : tone = `NM10;
		13'd155 : tone = `NM10;
		13'd156 : tone = `NM10;
		13'd157 : tone = `NM10;
		13'd158 : tone = `NM10;
		13'd159 : tone = `NM10;
		
		13'd160 : tone = `NM0;
		13'd161 : tone = `NM0;
		13'd162 : tone = `NM0;
		13'd163 : tone = `NM0;
		13'd164 : tone = `NM0;
		13'd165 : tone = `NM0;
		13'd166 : tone = `NM0;
		13'd167 : tone = `NM0;
		13'd168 : tone = `NM0;
		13'd169 : tone = `NM0;
		13'd170 : tone = `NM0;
		13'd171 : tone = `NM0;
		13'd172 : tone = `NM10;
		13'd173 : tone = `NM10;
		13'd174 : tone = `NM10;
		13'd175 : tone = `NM10;
		
		13'd176 : tone = `NM0;
		13'd177 : tone = `NM10;
		13'd178 : tone = `NM10;
		13'd179 : tone = `NM10;
		13'd180 : tone = `NM10;
		13'd181 : tone = `NM0;
		13'd182 : tone = `NM10;
		13'd183 : tone = `NM10;
		13'd184 : tone = `NM10;
		13'd185 : tone = `NM10;
		13'd186 : tone = `NM0;
		13'd187 : tone = `NM10;
		13'd188 : tone = `NM10;
		13'd189 : tone = `NM10;
		13'd190 : tone = `NM10;
		13'd191 : tone = `NM0;
		
		13'd192 : tone = `NM10;
		13'd193 : tone = `NM10;
		13'd194 : tone = `NM10;
		13'd195 : tone = `NM10;
		13'd196 : tone = `NM10;
		13'd197 : tone = `NM10;
		13'd198 : tone = `NM10;
		13'd199 : tone = `NM10;
		13'd200 : tone = `NM0;
		13'd201 : tone = `NM5;
		13'd202 : tone = `NM5;
		13'd203 : tone = `NM5;
		13'd204 : tone = `NM0;
		13'd205 : tone = `NM5;
		13'd206 : tone = `NM5;
		13'd207 : tone = `NM5;
		
		13'd208 : tone = `NM0;
		13'd209 : tone = `NM5;
		13'd210 : tone = `NM5;
		13'd211 : tone = `NM5;
		13'd212 : tone = `NM5;
		13'd213 : tone = `NM5;
		13'd214 : tone = `NM5;
		13'd215 : tone = `NM5;
		13'd216 : tone = `NM0;
		13'd217 : tone = `NM5;
		13'd218 : tone = `NM5;
		13'd219 : tone = `NM5;
		13'd220 : tone = `NM0;
		13'd221 : tone = `NM5;
		13'd222 : tone = `NM5;
		13'd223 : tone = `NM5;
		13'd224 : tone = `NM0;
		13'd225 : tone = `NM5;
		13'd226 : tone = `NM5;
		13'd227 : tone = `NM5;
		13'd228 : tone = `NM5;
		13'd229 : tone = `NM5;
		13'd230 : tone = `NM5;
		13'd231 : tone = `NM5;
		13'd232 : tone = `NM0;
		13'd233 : tone = `NM5;
		13'd234 : tone = `NM5;
		13'd235 : tone = `NM5;
		13'd236 : tone = `NM0;
		13'd237 : tone = `NM5;
		13'd238 : tone = `NM5;
		13'd239 : tone = `NM5;
		
		13'd240 : tone = `NM0;
		13'd241 : tone = `NM5;
		13'd242 : tone = `NM5;
		13'd243 : tone = `NM5;
		13'd244 : tone = `NM5;
		13'd245 : tone = `NM5;
		13'd246 : tone = `NM5;
		13'd247 : tone = `NM5;
		13'd248 : tone = `NM0;
		13'd249 : tone = `NM5;
		13'd250 : tone = `NM5;
		13'd251 : tone = `NM5;
		13'd252 : tone = `NM5;
		13'd253 : tone = `NM5;
		13'd254 : tone = `NM5;
		13'd255 : tone = `NM5;
		//repeat here
		13'd256: tone = `NM10;
        13'd257: tone = `NM10;
        13'd258: tone = `NM10;
        13'd259: tone = `NM10;
        13'd260: tone = `NM10;
        13'd261: tone = `NM10;
        13'd262: tone = `NM10;
        13'd263: tone = `NM10;
        13'd264: tone = `NM10;
        13'd265: tone = `NM10;
        13'd266: tone = `NM10;
        13'd267: tone = `NM10;
        13'd268: tone = `NM10;
        13'd269: tone = `NM10;
        13'd270: tone = `NM10;
        13'd271: tone = `NM0;
        
        13'd272: tone = `NM5;
        13'd273: tone = `NM5;
        13'd274: tone = `NM5;
        13'd275: tone = `NM5;
        13'd276: tone = `NM5;
        13'd277: tone = `NM5;
        13'd278: tone = `NM5;
        13'd279: tone = `NM5;
        13'd280: tone = `NM5;
        13'd281: tone = `NM5;
        13'd282: tone = `NM5;
        13'd283: tone = `NM5;
        13'd284: tone = `NM5;
        13'd285: tone = `NM5;
        13'd286: tone = `NM5;
        13'd287: tone = `NM5;
        
        13'd288: tone = `NM5;
        13'd289: tone = `NM5;
        13'd290: tone = `NM5;
        13'd291: tone = `NM5;
        13'd292: tone = `NM5;
        13'd293: tone = `NM5;
        13'd294: tone = `NM5;
        13'd295: tone = `NM0;
        13'd296: tone = `NM10;
        13'd297: tone = `NM10;
        13'd298: tone = `NM10;
        13'd299: tone = `NM10;
        13'd300: tone = `NM10;
        13'd301: tone = `NM10;
        13'd302: tone = `NM10;
        13'd303: tone = `NM0;
        
        13'd304: tone = `NM10;
        13'd305: tone = `NM10;
        13'd306: tone = `NM10;
        13'd307: tone = `NM10;
        13'd308: tone = `NM11;
        13'd309: tone = `NM11;
        13'd310: tone = `NM11;
        13'd311: tone = `NM11;
        13'd312: tone = `NM2 << 1; 
        13'd313: tone = `NM2 << 1;
        13'd314: tone = `NM2 << 1;
        13'd315: tone = `NM2 << 1;
        13'd316: tone = `NM3 << 1;
        13'd317: tone = `NM3 << 1;
        13'd318: tone = `NM3 << 1;
        13'd319: tone = `NM3 << 1;
        
        13'd320: tone = `NM5 << 1;
        13'd321: tone = `NM5 << 1;
        13'd322: tone = `NM5 << 1;
        13'd323: tone = `NM5 << 1;
        13'd324: tone = `NM5 << 1;
        13'd325: tone = `NM5 << 1;
        13'd326: tone = `NM5 << 1;
        13'd327: tone = `NM5 << 1;
        13'd328: tone = `NM5 << 1;
        13'd329: tone = `NM5 << 1;
        13'd330: tone = `NM5 << 1;
        13'd331: tone = `NM5 << 1;
        13'd332: tone = `NM5 << 1;
        13'd333: tone = `NM5 << 1;
        13'd334: tone = `NM5 << 1;
        13'd335: tone = `NM5 << 1;
        
        13'd336: tone = `NM5 << 1;
        13'd337: tone = `NM5 << 1;
        13'd338: tone = `NM5 << 1;
        13'd339: tone = `NM5 << 1;
        13'd340: tone = `NM5 << 1;
        13'd341: tone = `NM5 << 1;
        13'd342: tone = `NM5 << 1;
        13'd343: tone = `NM5 << 1;
        13'd344: tone = `NM5 << 1;
        13'd345: tone = `NM5 << 1;
        13'd346: tone = `NM5 << 1;
        13'd347: tone = `NM5 << 1;
        13'd348: tone = `NM5 << 1;
        13'd349: tone = `NM5 << 1;
        13'd350: tone = `NM5 << 1;
        13'd351: tone = `NM5 << 1;
        
        13'd352: tone = `NM0;
        13'd353: tone = `NM0;
        13'd354: tone = `NM0;
        13'd355: tone = `NM0;
        13'd356: tone = `NM0;
        13'd357: tone = `NM0;
        13'd358: tone = `NM0;
        13'd359: tone = `NM0;
        13'd360: tone = `NM5 << 1;
        13'd361: tone = `NM5 << 1;
        13'd362: tone = `NM5 << 1;
        13'd363: tone = `NM5 << 1;
        13'd364: tone = `NM5 << 1;
        13'd365: tone = `NM5 << 1;
        13'd366: tone = `NM5 << 1;
        13'd367: tone = `NM5 << 1;
        
        13'd368: tone = `NM0;
        13'd369: tone = `NM5 << 1;
        13'd370: tone = `NM5 << 1;
        13'd371: tone = `NM5 << 1;
        13'd372: tone = `NM5 << 1;
        13'd373: tone = `NM0;
        13'd374: tone = `NM6 << 1;
        13'd375: tone = `NM6 << 1;
        13'd376: tone = `NM6 << 1;
        13'd377: tone = `NM6 << 1;
        13'd378: tone = `NM0;
        13'd379: tone = `NM8 << 1;
        13'd380: tone = `NM8 << 1;
        13'd381: tone = `NM8 << 1;
        13'd382: tone = `NM8 << 1;
        13'd383: tone = `NM0;
        
        13'd384: tone = `NM10 << 1;
        13'd385: tone = `NM10 << 1;
        13'd386: tone = `NM10 << 1;
        13'd387: tone = `NM10 << 1;
        13'd388: tone = `NM10 << 1;
        13'd389: tone = `NM10 << 1;
        13'd390: tone = `NM10 << 1;
        13'd391: tone = `NM10 << 1;
        13'd392: tone = `NM10 << 1;
        13'd393: tone = `NM10 << 1;
        13'd394: tone = `NM10 << 1;
        13'd395: tone = `NM10 << 1;
        13'd396: tone = `NM10 << 1;
        13'd397: tone = `NM10 << 1;
        13'd398: tone = `NM10 << 1;
        13'd399: tone = `NM10 << 1;
        
        13'd400: tone = `NM10 << 1;
        13'd401: tone = `NM10 << 1;
        13'd402: tone = `NM10 << 1;
        13'd403: tone = `NM10 << 1;
        13'd404: tone = `NM10 << 1;
        13'd405: tone = `NM10 << 1;
        13'd406: tone = `NM10 << 1;
        13'd407: tone = `NM10 << 1;
        13'd408: tone = `NM10 << 1;
        13'd409: tone = `NM10 << 1;
        13'd410: tone = `NM10 << 1;
        13'd411: tone = `NM10 << 1;
        13'd412: tone = `NM10 << 1;
        13'd413: tone = `NM10 << 1;
        13'd414: tone = `NM10 << 1;
        13'd415: tone = `NM10 << 1;
        
        13'd416: tone = `NM0;
        13'd417: tone = `NM0;
        13'd418: tone = `NM0;
        13'd419: tone = `NM0;
        13'd420: tone = `NM0;
        13'd421: tone = `NM0;
        13'd422: tone = `NM0;
        13'd423: tone = `NM0;
        13'd424: tone = `NM10 << 1;
        13'd425: tone = `NM10 << 1;
        13'd426: tone = `NM10 << 1;
        13'd427: tone = `NM10 << 1;
        13'd428: tone = `NM10 << 1;
        13'd429: tone = `NM10 << 1;
        13'd430: tone = `NM10 << 1;
        13'd431: tone = `NM10 << 1;
        
        13'd432: tone = `NM0;
        13'd433: tone = `NM10 << 1;
        13'd434: tone = `NM10 << 1;
        13'd435: tone = `NM10 << 1;
        13'd436: tone = `NM10 << 1;
        13'd437: tone = `NM0;
        13'd438: tone = `NM8 << 1;
        13'd439: tone = `NM8 << 1;
        13'd440: tone = `NM8 << 1;
        13'd441: tone = `NM8 << 1;
        13'd442: tone = `NM0;
        13'd443: tone = `NM6 << 1;
        13'd444: tone = `NM6 << 1;
        13'd445: tone = `NM6 << 1;
        13'd446: tone = `NM6 << 1;
        13'd447: tone = `NM0;
        
        13'd448: tone = `NM8 << 1;
        13'd449: tone = `NM8 << 1;
        13'd450: tone = `NM8 << 1;
        13'd451: tone = `NM8 << 1;
        13'd452: tone = `NM8 << 1;
        13'd453: tone = `NM8 << 1;
        13'd454: tone = `NM8 << 1;
        13'd455: tone = `NM8 << 1;
        13'd456: tone = `NM8 << 1;
        13'd457: tone = `NM8 << 1;
        13'd458: tone = `NM8 << 1;
        13'd459: tone = `NM8 << 1;
        13'd460: tone = `NM6 << 1;
        13'd461: tone = `NM6 << 1;
        13'd462: tone = `NM6 << 1;
        13'd463: tone = `NM6 << 1;
        
        13'd464: tone = `NM5 << 1;
        13'd465: tone = `NM5 << 1;
        13'd466: tone = `NM5 << 1;
        13'd467: tone = `NM5 << 1;
        13'd468: tone = `NM5 << 1;
        13'd469: tone = `NM5 << 1;
        13'd470: tone = `NM5 << 1;
        13'd471: tone = `NM5 << 1;
        13'd472: tone = `NM5 << 1;
        13'd473: tone = `NM5 << 1;
        13'd474: tone = `NM5 << 1;
        13'd475: tone = `NM5 << 1;
        13'd476: tone = `NM5 << 1;
        13'd477: tone = `NM5 << 1;
        13'd478: tone = `NM5 << 1;
        13'd479: tone = `NM5 << 1;
        
        13'd480: tone = `NM5 << 1;
        13'd481: tone = `NM5 << 1;
        13'd482: tone = `NM5 << 1;
        13'd483: tone = `NM5 << 1;
        13'd484: tone = `NM5 << 1;
        13'd485: tone = `NM5 << 1;
        13'd486: tone = `NM5 << 1;
        13'd487: tone = `NM5 << 1;
        13'd488: tone = `NM5 << 1;
        13'd489: tone = `NM5 << 1;
        13'd490: tone = `NM5 << 1;
        13'd491: tone = `NM5 << 1;
        13'd492: tone = `NM5 << 1;
        13'd493: tone = `NM5 << 1;
        13'd494: tone = `NM5 << 1;
        13'd495: tone = `NM0;
        
        13'd496: tone = `NM5 << 1;
        13'd497: tone = `NM5 << 1;
        13'd498: tone = `NM5 << 1;
        13'd499: tone = `NM5 << 1;
        13'd500: tone = `NM5 << 1;
        13'd501: tone = `NM5 << 1;
        13'd502: tone = `NM5 << 1;
        13'd503: tone = `NM5 << 1;
        13'd504: tone = `NM5 << 1;
        13'd505: tone = `NM5 << 1;
        13'd506: tone = `NM5 << 1;
        13'd507: tone = `NM5 << 1;
        13'd508: tone = `NM5 << 1;
        13'd509: tone = `NM5 << 1;
        13'd510: tone = `NM5 << 1;
        13'd511: tone = `NM5 << 1;
        
        13'd512: tone = `NM3 << 1;
        13'd513: tone = `NM3 << 1;
        13'd514: tone = `NM3 << 1;
        13'd515: tone = `NM3 << 1;
        13'd516: tone = `NM3 << 1;
        13'd517: tone = `NM3 << 1;
        13'd518: tone = `NM3 << 1;
        13'd519: tone = `NM0;
        13'd520: tone = `NM3 << 1;
        13'd521: tone = `NM3 << 1;
        13'd522: tone = `NM3 << 1;
        13'd523: tone = `NM3 << 1;
        13'd524: tone = `NM5 << 1;
        13'd525: tone = `NM5 << 1;
        13'd526: tone = `NM5 << 1;
        13'd527: tone = `NM5 << 1;
        
        13'd528: tone = `NM6 << 1;
        13'd529: tone = `NM6 << 1;
        13'd530: tone = `NM6 << 1;
        13'd531: tone = `NM6 << 1;
        13'd532: tone = `NM6 << 1;
        13'd533: tone = `NM6 << 1;
        13'd534: tone = `NM6 << 1;
        13'd535: tone = `NM6 << 1;
        13'd536: tone = `NM6 << 1;
        13'd537: tone = `NM6 << 1;
        13'd538: tone = `NM6 << 1;
        13'd539: tone = `NM6 << 1;
        13'd540: tone = `NM6 << 1;
        13'd541: tone = `NM6 << 1;
        13'd542: tone = `NM6 << 1;
        13'd543: tone = `NM6 << 1;
        
        13'd544: tone = `NM6 << 1;
        13'd545: tone = `NM6 << 1;
        13'd546: tone = `NM6 << 1;
        13'd547: tone = `NM6 << 1;
        13'd548: tone = `NM6 << 1;
        13'd549: tone = `NM6 << 1;
        13'd550: tone = `NM6 << 1;
        13'd551: tone = `NM6 << 1;
        13'd552: tone = `NM6 << 1;
        13'd553: tone = `NM6 << 1;
        13'd554: tone = `NM6 << 1;
        13'd555: tone = `NM6 << 1;
        13'd556: tone = `NM6 << 1;
        13'd557: tone = `NM6 << 1;
        13'd558: tone = `NM6 << 1;
        13'd559: tone = `NM6 << 1;
        
        13'd560: tone = `NM5 << 1;
        13'd561: tone = `NM5 << 1;
        13'd562: tone = `NM5 << 1;
        13'd563: tone = `NM5 << 1;
        13'd564: tone = `NM5 << 1;
        13'd565: tone = `NM5 << 1;
        13'd566: tone = `NM5 << 1;
        13'd567: tone = `NM5 << 1;
        13'd568: tone = `NM3 << 1;
        13'd569: tone = `NM3 << 1;
        13'd570: tone = `NM3 << 1;
        13'd571: tone = `NM3 << 1;
        13'd572: tone = `NM3 << 1;
        13'd573: tone = `NM3 << 1;
        13'd574: tone = `NM3 << 1;
        13'd575: tone = `NM3 << 1;
        
        13'd576: tone = `NM1 << 1;
        13'd577: tone = `NM1 << 1;
        13'd578: tone = `NM1 << 1;
        13'd579: tone = `NM1 << 1;
        13'd580: tone = `NM1 << 1;
        13'd581: tone = `NM1 << 1;
        13'd582: tone = `NM1 << 1;
        13'd583: tone = `NM0;
        13'd584: tone = `NM1 << 1;
        13'd585: tone = `NM1 << 1;
        13'd586: tone = `NM1 << 1;
        13'd587: tone = `NM1 << 1;
        13'd588: tone = `NM3 << 1;
        13'd589: tone = `NM3 << 1;
        13'd590: tone = `NM3 << 1;
        13'd591: tone = `NM3 << 1;
        
        13'd592: tone = `NM5 << 1;
        13'd593: tone = `NM5 << 1;
        13'd594: tone = `NM5 << 1;
        13'd595: tone = `NM5 << 1;
        13'd596: tone = `NM5 << 1;
        13'd597: tone = `NM5 << 1;
        13'd598: tone = `NM5 << 1;
        13'd599: tone = `NM5 << 1;
        13'd600: tone = `NM5 << 1;
        13'd601: tone = `NM5 << 1;
        13'd602: tone = `NM5 << 1;
        13'd603: tone = `NM5 << 1;
        13'd604: tone = `NM5 << 1;
        13'd605: tone = `NM5 << 1;
        13'd606: tone = `NM5 << 1;
        13'd607: tone = `NM5 << 1;
        
        13'd608: tone = `NM5 << 1;
        13'd609: tone = `NM5 << 1;
        13'd610: tone = `NM5 << 1;
        13'd611: tone = `NM5 << 1;
        13'd612: tone = `NM5 << 1;
        13'd613: tone = `NM5 << 1;
        13'd614: tone = `NM5 << 1;
        13'd615: tone = `NM5 << 1;
        13'd616: tone = `NM5 << 1;
        13'd617: tone = `NM5 << 1;
        13'd618: tone = `NM5 << 1;
        13'd619: tone = `NM5 << 1;
        13'd620: tone = `NM5 << 1;
        13'd621: tone = `NM5 << 1;
        13'd622: tone = `NM5 << 1;
        13'd623: tone = `NM5 << 1;
        
        13'd624: tone = `NM3 << 1;
        13'd625: tone = `NM3 << 1;
        13'd626: tone = `NM3 << 1;
        13'd627: tone = `NM3 << 1;
        13'd628: tone = `NM3 << 1;
        13'd629: tone = `NM3 << 1;
        13'd630: tone = `NM3 << 1;
        13'd631: tone = `NM3 << 1;
        13'd632: tone = `NM1 << 1;
        13'd633: tone = `NM1 << 1;
        13'd634: tone = `NM1 << 1;
        13'd635: tone = `NM1 << 1;
        13'd636: tone = `NM1 << 1;
        13'd637: tone = `NM1 << 1;
        13'd638: tone = `NM1 << 1;
        13'd639: tone = `NM1 << 1;
        
        13'd640: tone = `NM11;
        13'd641: tone = `NM11;
        13'd642: tone = `NM11;
        13'd643: tone = `NM11;
        13'd644: tone = `NM11;
        13'd645: tone = `NM11;
        13'd646: tone = `NM11;
        13'd647: tone = `NM0;
        13'd648: tone = `NM11;
        13'd649: tone = `NM11;
        13'd650: tone = `NM11;
        13'd651: tone = `NM11;
        13'd652: tone = `NM2 << 1;
        13'd653: tone = `NM2 << 1;
        13'd654: tone = `NM2 << 1;
        13'd655: tone = `NM2 << 1;
        
        13'd656: tone = `NM4 << 1;
        13'd657: tone = `NM4 << 1;
        13'd658: tone = `NM4 << 1;
        13'd659: tone = `NM4 << 1;
        13'd660: tone = `NM4 << 1;
        13'd661: tone = `NM4 << 1;
        13'd662: tone = `NM4 << 1;
        13'd663: tone = `NM4 << 1;
        13'd664: tone = `NM4 << 1;
        13'd665: tone = `NM4 << 1;
        13'd666: tone = `NM4 << 1;
        13'd667: tone = `NM4 << 1;
        13'd668: tone = `NM4 << 1;
        13'd669: tone = `NM4 << 1;
        13'd670: tone = `NM4 << 1;
        13'd671: tone = `NM4 << 1;
        
        13'd672: tone = `NM4 << 1;
        13'd673: tone = `NM4 << 1;
        13'd674: tone = `NM4 << 1;
        13'd675: tone = `NM4 << 1;
        13'd676: tone = `NM4 << 1;
        13'd677: tone = `NM4 << 1;
        13'd678: tone = `NM4 << 1;
        13'd679: tone = `NM4 << 1;
        13'd680: tone = `NM4 << 1;
        13'd681: tone = `NM4 << 1;
        13'd682: tone = `NM4 << 1;
        13'd683: tone = `NM4 << 1;
        13'd684: tone = `NM4 << 1;
        13'd685: tone = `NM4 << 1;
        13'd686: tone = `NM4 << 1;
        13'd687: tone = `NM4 << 1;
        
        13'd688: tone = `NM7 << 1;
        13'd689: tone = `NM7 << 1;
        13'd690: tone = `NM7 << 1;
        13'd691: tone = `NM7 << 1;
        13'd692: tone = `NM7 << 1;
        13'd693: tone = `NM7 << 1;
        13'd694: tone = `NM7 << 1;
        13'd695: tone = `NM7 << 1;
        13'd696: tone = `NM7 << 1;
        13'd697: tone = `NM7 << 1;
        13'd698: tone = `NM7 << 1;
        13'd699: tone = `NM7 << 1;
        13'd700: tone = `NM7 << 1;
        13'd701: tone = `NM7 << 1;
        13'd702: tone = `NM7 << 1;
        13'd703: tone = `NM7 << 1;
        
        13'd704: tone = `NM5 << 1;
        13'd705: tone = `NM5 << 1;
        13'd706: tone = `NM5 << 1;
        13'd707: tone = `NM5 << 1;
        13'd708: tone = `NM5 << 1;
        13'd709: tone = `NM5 << 1;
        13'd710: tone = `NM5 << 1;
        13'd711: tone = `NM5 << 1;
        13'd712: tone = `NM5;
        13'd713: tone = `NM5;
        13'd714: tone = `NM5;
        13'd715: tone = `NM0;
        13'd716: tone = `NM5;
        13'd717: tone = `NM5;
        13'd718: tone = `NM5;
        13'd719: tone = `NM0;
        
        13'd720: tone = `NM5;
        13'd721: tone = `NM5;
        13'd722: tone = `NM5;
        13'd723: tone = `NM5;
        13'd724: tone = `NM5;
        13'd725: tone = `NM5;
        13'd726: tone = `NM5;
        13'd727: tone = `NM0;
        13'd728: tone = `NM5;
        13'd729: tone = `NM5;
        13'd730: tone = `NM5;
        13'd731: tone = `NM0;
        13'd732: tone = `NM5;
        13'd733: tone = `NM5;
        13'd734: tone = `NM5;
        13'd735: tone = `NM0;
        
        13'd736: tone = `NM5;
        13'd737: tone = `NM5;
        13'd738: tone = `NM5;
        13'd739: tone = `NM5;
        13'd740: tone = `NM5;
        13'd741: tone = `NM5;
        13'd742: tone = `NM5;
        13'd743: tone = `NM0;
        13'd744: tone = `NM5;
        13'd745: tone = `NM5;
        13'd746: tone = `NM5;
        13'd747: tone = `NM0;
        13'd748: tone = `NM5;
        13'd749: tone = `NM5;
        13'd750: tone = `NM5;
        13'd751: tone = `NM0;
        
        13'd752: tone = `NM5;
        13'd753: tone = `NM5;
        13'd754: tone = `NM5;
        13'd755: tone = `NM5;
        13'd756: tone = `NM5;
        13'd757: tone = `NM5;
        13'd758: tone = `NM5;
        13'd759: tone = `NM0;
        13'd760: tone = `NM5;
        13'd761: tone = `NM5;
        13'd762: tone = `NM5;
        13'd763: tone = `NM5;
        13'd764: tone = `NM5;
        13'd765: tone = `NM5;
        13'd766: tone = `NM5;
        13'd767: tone = `NM5;
        
        13'd768: tone = `NM10;
        13'd769: tone = `NM10;
        13'd770: tone = `NM10;
        13'd771: tone = `NM10;
        13'd772: tone = `NM10;
        13'd773: tone = `NM10;
        13'd774: tone = `NM10;
        13'd775: tone = `NM10;
        13'd776: tone = `NM10;
        13'd777: tone = `NM10;
        13'd778: tone = `NM10;
        13'd779: tone = `NM10;
        13'd780: tone = `NM10;
        13'd781: tone = `NM10;
        13'd782: tone = `NM10;
        13'd783: tone = `NM10;
        
        13'd784: tone = `NM5;
        13'd785: tone = `NM5;
        13'd786: tone = `NM5;
        13'd787: tone = `NM5;
        13'd788: tone = `NM5;
        13'd789: tone = `NM5;
        13'd790: tone = `NM5;
        13'd791: tone = `NM5;
        13'd792: tone = `NM5;
        13'd793: tone = `NM5;
        13'd794: tone = `NM5;
        13'd795: tone = `NM5;
        13'd796: tone = `NM5;
        13'd797: tone = `NM5;
        13'd798: tone = `NM5;
        13'd799: tone = `NM5;
        
        13'd800: tone = `NM5;
        13'd801: tone = `NM5;
        13'd802: tone = `NM5;
        13'd803: tone = `NM5;
        13'd804: tone = `NM5;
        13'd805: tone = `NM5;
        13'd806: tone = `NM5;
        13'd807: tone = `NM5;
        13'd808: tone = `NM10;
        13'd809: tone = `NM10;
        13'd810: tone = `NM10;
        13'd811: tone = `NM10;
        13'd812: tone = `NM10;
        13'd813: tone = `NM10;
        13'd814: tone = `NM10;
        13'd815: tone = `NM0;
        
        13'd816: tone = `NM10;
        13'd817: tone = `NM10;
        13'd818: tone = `NM10;
        13'd819: tone = `NM10;
        13'd820: tone = `NM11;
        13'd821: tone = `NM11;
        13'd822: tone = `NM11;
        13'd823: tone = `NM11;
        13'd824: tone = `NM2 << 1;
        13'd825: tone = `NM2 << 1;
        13'd826: tone = `NM2 << 1;
        13'd827: tone = `NM2 << 1;
        13'd828: tone = `NM3 << 1;
        13'd829: tone = `NM3 << 1;
        13'd830: tone = `NM3 << 1;
        13'd831: tone = `NM3 << 1;
        
        13'd832: tone = `NM5 << 1;
        13'd833: tone = `NM5 << 1;
        13'd834: tone = `NM5 << 1;
        13'd835: tone = `NM5 << 1;
        13'd836: tone = `NM5 << 1;
        13'd837: tone = `NM5 << 1;
        13'd838: tone = `NM5 << 1;
        13'd839: tone = `NM5 << 1;
        13'd840: tone = `NM5 << 1;
        13'd841: tone = `NM5 << 1;
        13'd842: tone = `NM5 << 1;
        13'd843: tone = `NM5 << 1;
        13'd844: tone = `NM5 << 1;
        13'd845: tone = `NM5 << 1;
        13'd846: tone = `NM5 << 1;
        13'd847: tone = `NM5 << 1;
        
        13'd848: tone = `NM5 << 1;
        13'd849: tone = `NM5 << 1;
        13'd850: tone = `NM5 << 1;
        13'd851: tone = `NM5 << 1;
        13'd852: tone = `NM5 << 1;
        13'd853: tone = `NM5 << 1;
        13'd854: tone = `NM5 << 1;
        13'd855: tone = `NM5 << 1;
        13'd856: tone = `NM5 << 1;
        13'd857: tone = `NM5 << 1;
        13'd858: tone = `NM5 << 1;
        13'd859: tone = `NM5 << 1;
        13'd860: tone = `NM5 << 1;
        13'd861: tone = `NM5 << 1;
        13'd862: tone = `NM5 << 1;
        13'd863: tone = `NM5 << 1;
        
        13'd864: tone = `NM0;
        13'd865: tone = `NM0;
        13'd866: tone = `NM0;
        13'd867: tone = `NM0;
        13'd868: tone = `NM0;
        13'd869: tone = `NM0;
        13'd870: tone = `NM0;
        13'd871: tone = `NM0;
        13'd872: tone = `NM5 << 1;
        13'd873: tone = `NM5 << 1;
        13'd874: tone = `NM5 << 1;
        13'd875: tone = `NM5 << 1;
        13'd876: tone = `NM5 << 1;
        13'd877: tone = `NM5 << 1;
        13'd878: tone = `NM5 << 1;
        13'd879: tone = `NM5 << 1;
        
        13'd880: tone = `NM0;
        13'd881: tone = `NM5 << 1;
        13'd882: tone = `NM5 << 1;
        13'd883: tone = `NM5 << 1;
        13'd884: tone = `NM5 << 1;
        13'd885: tone = `NM0;
        13'd886: tone = `NM6 << 1;
        13'd887: tone = `NM6 << 1;
        13'd888: tone = `NM6 << 1;
        13'd889: tone = `NM6 << 1;
        13'd890: tone = `NM0;
        13'd891: tone = `NM8 << 1;
        13'd892: tone = `NM8 << 1;
        13'd893: tone = `NM8 << 1;
        13'd894: tone = `NM8 << 1;
        13'd895: tone = `NM0;
        
        13'd896: tone = `NM10 << 1;
        13'd897: tone = `NM10 << 1;
        13'd898: tone = `NM10 << 1;
        13'd899: tone = `NM10 << 1;
        13'd900: tone = `NM10 << 1;
        13'd901: tone = `NM10 << 1;
        13'd902: tone = `NM10 << 1;
        13'd903: tone = `NM10 << 1;
        13'd904: tone = `NM10 << 1;
        13'd905: tone = `NM10 << 1;
        13'd906: tone = `NM10 << 1;
        13'd907: tone = `NM10 << 1;
        13'd908: tone = `NM10 << 1;
        13'd909: tone = `NM10 << 1;
        13'd910: tone = `NM10 << 1;
        13'd911: tone = `NM10 << 1;
        
        13'd912: tone = `NM0;
        13'd913: tone = `NM0;
        13'd914: tone = `NM0;
        13'd915: tone = `NM0;
        13'd916: tone = `NM0;
        13'd917: tone = `NM0;
        13'd918: tone = `NM0;
        13'd919: tone = `NM0;
        13'd920: tone = `NM0;
        13'd921: tone = `NM0;
        13'd922: tone = `NM0;
        13'd923: tone = `NM0;
        13'd924: tone = `NM0;
        13'd925: tone = `NM0;
        13'd926: tone = `NM0;
        13'd927: tone = `NM0;
        
        13'd928: tone = `NM1 << 2;
        13'd929: tone = `NM1 << 2;
        13'd930: tone = `NM1 << 2;
        13'd931: tone = `NM1 << 2;
        13'd932: tone = `NM1 << 2;
        13'd933: tone = `NM1 << 2;
        13'd934: tone = `NM1 << 2;
        13'd935: tone = `NM1 << 2;
        13'd936: tone = `NM1 << 2;
        13'd937: tone = `NM1 << 2;
        13'd938: tone = `NM1 << 2;
        13'd939: tone = `NM1 << 2;
        13'd940: tone = `NM1 << 2;
        13'd941: tone = `NM1 << 2;
        13'd942: tone = `NM1 << 2;
        13'd943: tone = `NM1 << 2;
        
        13'd944: tone = `NM11 << 1;
        13'd945: tone = `NM11 << 1;
        13'd946: tone = `NM11 << 1;
        13'd947: tone = `NM11 << 1;
        13'd948: tone = `NM11 << 1;
        13'd949: tone = `NM11 << 1;
        13'd950: tone = `NM11 << 1;
        13'd951: tone = `NM11 << 1;
        13'd952: tone = `NM11 << 1;
        13'd953: tone = `NM11 << 1;
        13'd954: tone = `NM11 << 1;
        13'd955: tone = `NM11 << 1;
        13'd956: tone = `NM11 << 1;
        13'd957: tone = `NM11 << 1;
        13'd958: tone = `NM11 << 1;
        13'd959: tone = `NM11 << 1;
        
        13'd960: tone = `NM9 << 1;
        13'd961: tone = `NM9 << 1;
        13'd962: tone = `NM9 << 1;
        13'd963: tone = `NM9 << 1;
        13'd964: tone = `NM9 << 1;
        13'd965: tone = `NM9 << 1;
        13'd966: tone = `NM9 << 1;
        13'd967: tone = `NM9 << 1;
        13'd968: tone = `NM9 << 1;
        13'd969: tone = `NM9 << 1;
        13'd970: tone = `NM9 << 1;
        13'd971: tone = `NM9 << 1;
        13'd972: tone = `NM9 << 1;
        13'd973: tone = `NM9 << 1;
        13'd974: tone = `NM9 << 1;
        13'd975: tone = `NM9 << 1;
        
        13'd976: tone = `NM9 << 1;
        13'd977: tone = `NM9 << 1;
        13'd978: tone = `NM9 << 1;
        13'd979: tone = `NM9 << 1;
        13'd980: tone = `NM9 << 1;
        13'd981: tone = `NM9 << 1;
        13'd982: tone = `NM9 << 1;
        13'd983: tone = `NM9 << 1;
        13'd984: tone = `NM9 << 1;
        13'd985: tone = `NM9 << 1;
        13'd986: tone = `NM9 << 1;
        13'd987: tone = `NM9 << 1;
        13'd988: tone = `NM9 << 1;
        13'd989: tone = `NM9 << 1;
        13'd990: tone = `NM9 << 1;
        13'd991: tone = `NM9 << 1;
        
        13'd992: tone = `NM5 << 1;
        13'd993: tone = `NM5 << 1;
        13'd994: tone = `NM5 << 1;
        13'd995: tone = `NM5 << 1;
        13'd996: tone = `NM5 << 1;
        13'd997: tone = `NM5 << 1;
        13'd998: tone = `NM5 << 1;
        13'd999: tone = `NM5 << 1;
        13'd1000: tone = `NM5 << 1;
        13'd1001: tone = `NM5 << 1;
        13'd1002: tone = `NM5 << 1;
        13'd1003: tone = `NM5 << 1;
        13'd1004: tone = `NM5 << 1;
        13'd1005: tone = `NM5 << 1;
        13'd1006: tone = `NM5 << 1;
        13'd1007: tone = `NM5 << 1;
        
        13'd1008: tone = `NM6 << 1;
        13'd1009: tone = `NM6 << 1;
        13'd1010: tone = `NM6 << 1;
        13'd1011: tone = `NM6 << 1;
        13'd1012: tone = `NM6 << 1;
        13'd1013: tone = `NM6 << 1;
        13'd1014: tone = `NM6 << 1;
        13'd1015: tone = `NM6 << 1;
        13'd1016: tone = `NM6 << 1;
        13'd1017: tone = `NM6 << 1;
        13'd1018: tone = `NM6 << 1;
        13'd1019: tone = `NM6 << 1;
        13'd1020: tone = `NM6 << 1;
        13'd1021: tone = `NM6 << 1;
        13'd1022: tone = `NM6 << 1;
        13'd1023: tone = `NM6 << 1;
        
        13'd1024: tone = `NM6 << 1;
        13'd1025: tone = `NM6 << 1;
        13'd1026: tone = `NM6 << 1;
        13'd1027: tone = `NM6 << 1;
        13'd1028: tone = `NM6 << 1;
        13'd1029: tone = `NM6 << 1;
        13'd1030: tone = `NM6 << 1;
        13'd1031: tone = `NM6 << 1;
        13'd1032: tone = `NM6 << 1;
        13'd1033: tone = `NM6 << 1;
        13'd1034: tone = `NM6 << 1;
        13'd1035: tone = `NM6 << 1;
        13'd1036: tone = `NM6 << 1;
        13'd1037: tone = `NM6 << 1;
        13'd1038: tone = `NM6 << 1;
        13'd1039: tone = `NM6 << 1;
        
        13'd1040: tone = `NM6 << 1;
        13'd1041: tone = `NM6 << 1;
        13'd1042: tone = `NM6 << 1;
        13'd1043: tone = `NM6 << 1;
        13'd1044: tone = `NM6 << 1;
        13'd1045: tone = `NM6 << 1;
        13'd1046: tone = `NM6 << 1;
        13'd1047: tone = `NM6 << 1;
        13'd1048: tone = `NM6 << 1;
        13'd1049: tone = `NM6 << 1;
        13'd1050: tone = `NM6 << 1;
        13'd1051: tone = `NM6 << 1;
        13'd1052: tone = `NM6 << 1;
        13'd1053: tone = `NM6 << 1;
        13'd1054: tone = `NM6 << 1;
        13'd1055: tone = `NM6 << 1;
        
        13'd1056: tone = `NM10 << 1;
        13'd1057: tone = `NM10 << 1;
        13'd1058: tone = `NM10 << 1;
        13'd1059: tone = `NM10 << 1;
        13'd1060: tone = `NM10 << 1;
        13'd1061: tone = `NM10 << 1;
        13'd1062: tone = `NM10 << 1;
        13'd1063: tone = `NM10 << 1;
        13'd1064: tone = `NM10 << 1;
        13'd1065: tone = `NM10 << 1;
        13'd1066: tone = `NM10 << 1;
        13'd1067: tone = `NM10 << 1;
        13'd1068: tone = `NM10 << 1;
        13'd1069: tone = `NM10 << 1;
        13'd1070: tone = `NM10 << 1;
        13'd1071: tone = `NM10 << 1;
        
        13'd1072: tone = `NM9 << 1;
        13'd1073: tone = `NM9 << 1;
        13'd1074: tone = `NM9 << 1;
        13'd1075: tone = `NM9 << 1;
        13'd1076: tone = `NM9 << 1;
        13'd1077: tone = `NM9 << 1;
        13'd1078: tone = `NM9 << 1;
        13'd1079: tone = `NM9 << 1;
        13'd1080: tone = `NM9 << 1;
        13'd1081: tone = `NM9 << 1;
        13'd1082: tone = `NM9 << 1;
        13'd1083: tone = `NM9 << 1;
        13'd1084: tone = `NM9 << 1;
        13'd1085: tone = `NM9 << 1;
        13'd1086: tone = `NM9 << 1;
        13'd1087: tone = `NM9 << 1;
        
        13'd1088: tone = `NM5 << 1;
        13'd1089: tone = `NM5 << 1;
        13'd1090: tone = `NM5 << 1;
        13'd1091: tone = `NM5 << 1;
        13'd1092: tone = `NM5 << 1;
        13'd1093: tone = `NM5 << 1;
        13'd1094: tone = `NM5 << 1;
        13'd1095: tone = `NM5 << 1;
        13'd1096: tone = `NM5 << 1;
        13'd1097: tone = `NM5 << 1;
        13'd1098: tone = `NM5 << 1;
        13'd1099: tone = `NM5 << 1;
        13'd1100: tone = `NM5 << 1;
        13'd1101: tone = `NM5 << 1;
        13'd1102: tone = `NM5 << 1;
        13'd1103: tone = `NM5 << 1;
        
        13'd1104: tone = `NM5 << 1;
        13'd1105: tone = `NM5 << 1;
        13'd1106: tone = `NM5 << 1;
        13'd1107: tone = `NM5 << 1;
        13'd1108: tone = `NM5 << 1;
        13'd1109: tone = `NM5 << 1;
        13'd1110: tone = `NM5 << 1;
        13'd1111: tone = `NM5 << 1;
        13'd1112: tone = `NM5 << 1;
        13'd1113: tone = `NM5 << 1;
        13'd1114: tone = `NM5 << 1;
        13'd1115: tone = `NM5 << 1;
        13'd1116: tone = `NM5 << 1;
        13'd1117: tone = `NM5 << 1;
        13'd1118: tone = `NM5 << 1;
        13'd1119: tone = `NM0;
        
        13'd1120: tone = `NM5 << 1;
        13'd1121: tone = `NM5 << 1;
        13'd1122: tone = `NM5 << 1;
        13'd1123: tone = `NM5 << 1;
        13'd1124: tone = `NM5 << 1;
        13'd1125: tone = `NM5 << 1;
        13'd1126: tone = `NM5 << 1;
        13'd1127: tone = `NM5 << 1;
        13'd1128: tone = `NM5 << 1;
        13'd1129: tone = `NM5 << 1;
        13'd1130: tone = `NM5 << 1;
        13'd1131: tone = `NM5 << 1;
        13'd1132: tone = `NM5 << 1;
        13'd1133: tone = `NM5 << 1;
        13'd1134: tone = `NM5 << 1;
        13'd1135: tone = `NM5 << 1;
        
        13'd1136: tone = `NM6 << 1;
        13'd1137: tone = `NM6 << 1;
        13'd1138: tone = `NM6 << 1;
        13'd1139: tone = `NM6 << 1;
        13'd1140: tone = `NM6 << 1;
        13'd1141: tone = `NM6 << 1;
        13'd1142: tone = `NM6 << 1;
        13'd1143: tone = `NM6 << 1;
        13'd1144: tone = `NM6 << 1;
        13'd1145: tone = `NM6 << 1;
        13'd1146: tone = `NM6 << 1;
        13'd1147: tone = `NM6 << 1;
        13'd1148: tone = `NM6 << 1;
        13'd1149: tone = `NM6 << 1;
        13'd1150: tone = `NM6 << 1;
        13'd1151: tone = `NM6 << 1;
        
        13'd1152: tone = `NM6 << 1;
        13'd1153: tone = `NM6 << 1;
        13'd1154: tone = `NM6 << 1;
        13'd1155: tone = `NM6 << 1;
        13'd1156: tone = `NM6 << 1;
        13'd1157: tone = `NM6 << 1;
        13'd1158: tone = `NM6 << 1;
        13'd1159: tone = `NM6 << 1;
        13'd1160: tone = `NM6 << 1;
        13'd1161: tone = `NM6 << 1;
        13'd1162: tone = `NM6 << 1;
        13'd1163: tone = `NM6 << 1;
        13'd1164: tone = `NM6 << 1;
        13'd1165: tone = `NM6 << 1;
        13'd1166: tone = `NM6 << 1;
        13'd1167: tone = `NM6 << 1;
        
        13'd1168: tone = `NM6 << 1;
        13'd1169: tone = `NM6 << 1;
        13'd1170: tone = `NM6 << 1;
        13'd1171: tone = `NM6 << 1;
        13'd1172: tone = `NM6 << 1;
        13'd1173: tone = `NM6 << 1;
        13'd1174: tone = `NM6 << 1;
        13'd1175: tone = `NM6 << 1;
        13'd1176: tone = `NM6 << 1;
        13'd1177: tone = `NM6 << 1;
        13'd1178: tone = `NM6 << 1;
        13'd1179: tone = `NM6 << 1;
        13'd1180: tone = `NM6 << 1;
        13'd1181: tone = `NM6 << 1;
        13'd1182: tone = `NM6 << 1;
        13'd1183: tone = `NM6 << 1;
        
        13'd1184: tone = `NM10 << 1;
        13'd1185: tone = `NM10 << 1;
        13'd1186: tone = `NM10 << 1;
        13'd1187: tone = `NM10 << 1;
        13'd1188: tone = `NM10 << 1;
        13'd1189: tone = `NM10 << 1;
        13'd1190: tone = `NM10 << 1;
        13'd1191: tone = `NM10 << 1;
        13'd1192: tone = `NM10 << 1;
        13'd1193: tone = `NM10 << 1;
        13'd1194: tone = `NM10 << 1;
        13'd1195: tone = `NM10 << 1;
        13'd1196: tone = `NM10 << 1;
        13'd1197: tone = `NM10 << 1;
        13'd1198: tone = `NM10 << 1;
        13'd1199: tone = `NM10 << 1;
        
        13'd1200: tone = `NM9 << 1;
        13'd1201: tone = `NM9 << 1;
        13'd1202: tone = `NM9 << 1;
        13'd1203: tone = `NM9 << 1;
        13'd1204: tone = `NM9 << 1;
        13'd1205: tone = `NM9 << 1;
        13'd1206: tone = `NM9 << 1;
        13'd1207: tone = `NM9 << 1;
        13'd1208: tone = `NM9 << 1;
        13'd1209: tone = `NM9 << 1;
        13'd1210: tone = `NM9 << 1;
        13'd1211: tone = `NM9 << 1;
        13'd1212: tone = `NM9 << 1;
        13'd1213: tone = `NM9 << 1;
        13'd1214: tone = `NM9 << 1;
        13'd1215: tone = `NM9 << 1;
        
        13'd1216: tone = `NM5 << 1;
        13'd1217: tone = `NM5 << 1;
        13'd1218: tone = `NM5 << 1;
        13'd1219: tone = `NM5 << 1;
        13'd1220: tone = `NM5 << 1;
        13'd1221: tone = `NM5 << 1;
        13'd1222: tone = `NM5 << 1;
        13'd1223: tone = `NM5 << 1;
        13'd1224: tone = `NM5 << 1;
        13'd1225: tone = `NM5 << 1;
        13'd1226: tone = `NM5 << 1;
        13'd1227: tone = `NM5 << 1;
        13'd1228: tone = `NM5 << 1;
        13'd1229: tone = `NM5 << 1;
        13'd1230: tone = `NM5 << 1;
        13'd1231: tone = `NM5 << 1;
        
        13'd1232: tone = `NM5 << 1;
        13'd1233: tone = `NM5 << 1;
        13'd1234: tone = `NM5 << 1;
        13'd1235: tone = `NM5 << 1;
        13'd1236: tone = `NM5 << 1;
        13'd1237: tone = `NM5 << 1;
        13'd1238: tone = `NM5 << 1;
        13'd1239: tone = `NM5 << 1;
        13'd1240: tone = `NM5 << 1;
        13'd1241: tone = `NM5 << 1;
        13'd1242: tone = `NM5 << 1;
        13'd1243: tone = `NM5 << 1;
        13'd1244: tone = `NM5 << 1;
        13'd1245: tone = `NM5 << 1;
        13'd1246: tone = `NM5 << 1;
        13'd1247: tone = `NM5 << 1;
        
        13'd1248: tone = `NM2 << 1;
        13'd1249: tone = `NM2 << 1;
        13'd1250: tone = `NM2 << 1;
        13'd1251: tone = `NM2 << 1;
        13'd1252: tone = `NM2 << 1;
        13'd1253: tone = `NM2 << 1;
        13'd1254: tone = `NM2 << 1;
        13'd1255: tone = `NM2 << 1;
        13'd1256: tone = `NM2 << 1;
        13'd1257: tone = `NM2 << 1;
        13'd1258: tone = `NM2 << 1;
        13'd1259: tone = `NM2 << 1;
        13'd1260: tone = `NM2 << 1;
        13'd1261: tone = `NM2 << 1;
        13'd1262: tone = `NM2 << 1;
        13'd1263: tone = `NM2 << 1;
        
        13'd1264: tone = `NM3 << 1;
        13'd1265: tone = `NM3 << 1;
        13'd1266: tone = `NM3 << 1;
        13'd1267: tone = `NM3 << 1;
        13'd1268: tone = `NM3 << 1;
        13'd1269: tone = `NM3 << 1;
        13'd1270: tone = `NM3 << 1;
        13'd1271: tone = `NM3 << 1;
        13'd1272: tone = `NM3 << 1;
        13'd1273: tone = `NM3 << 1;
        13'd1274: tone = `NM3 << 1;
        13'd1275: tone = `NM3 << 1;
        13'd1276: tone = `NM3 << 1;
        13'd1277: tone = `NM3 << 1;
        13'd1278: tone = `NM3 << 1;
        13'd1279: tone = `NM3 << 1;
        
        13'd1280: tone = `NM3 << 1;
        13'd1281: tone = `NM3 << 1;
        13'd1282: tone = `NM3 << 1;
        13'd1283: tone = `NM3 << 1;
        13'd1284: tone = `NM3 << 1;
        13'd1285: tone = `NM3 << 1;
        13'd1286: tone = `NM3 << 1;
        13'd1287: tone = `NM3 << 1;
        13'd1288: tone = `NM3 << 1;
        13'd1289: tone = `NM3 << 1;
        13'd1290: tone = `NM3 << 1;
        13'd1291: tone = `NM3 << 1;
        13'd1292: tone = `NM3 << 1;
        13'd1293: tone = `NM3 << 1;
        13'd1294: tone = `NM3 << 1;
        13'd1295: tone = `NM3 << 1;
        
        13'd1296: tone = `NM3 << 1;
        13'd1297: tone = `NM3 << 1;
        13'd1298: tone = `NM3 << 1;
        13'd1299: tone = `NM3 << 1;
        13'd1300: tone = `NM3 << 1;
        13'd1301: tone = `NM3 << 1;
        13'd1302: tone = `NM3 << 1;
        13'd1303: tone = `NM3 << 1;
        13'd1304: tone = `NM3 << 1;
        13'd1305: tone = `NM3 << 1;
        13'd1306: tone = `NM3 << 1;
        13'd1307: tone = `NM3 << 1;
        13'd1308: tone = `NM3 << 1;
        13'd1309: tone = `NM3 << 1;
        13'd1310: tone = `NM3 << 1;
        13'd1311: tone = `NM3 << 1;
        
        13'd1312: tone = `NM6 << 1;
        13'd1313: tone = `NM6 << 1;
        13'd1314: tone = `NM6 << 1;
        13'd1315: tone = `NM6 << 1;
        13'd1316: tone = `NM6 << 1;
        13'd1317: tone = `NM6 << 1;
        13'd1318: tone = `NM6 << 1;
        13'd1319: tone = `NM6 << 1;
        13'd1320: tone = `NM6 << 1;
        13'd1321: tone = `NM6 << 1;
        13'd1322: tone = `NM6 << 1;
        13'd1323: tone = `NM6 << 1;
        13'd1324: tone = `NM6 << 1;
        13'd1325: tone = `NM6 << 1;
        13'd1326: tone = `NM6 << 1;
        13'd1327: tone = `NM6 << 1;
        
        13'd1328: tone = `NM5 << 1;
        13'd1329: tone = `NM5 << 1;
        13'd1330: tone = `NM5 << 1;
        13'd1331: tone = `NM5 << 1;
        13'd1332: tone = `NM5 << 1;
        13'd1333: tone = `NM5 << 1;
        13'd1334: tone = `NM5 << 1;
        13'd1335: tone = `NM5 << 1;
        13'd1336: tone = `NM5 << 1;
        13'd1337: tone = `NM5 << 1;
        13'd1338: tone = `NM5 << 1;
        13'd1339: tone = `NM5 << 1;
        13'd1340: tone = `NM5 << 1;
        13'd1341: tone = `NM5 << 1;
        13'd1342: tone = `NM5 << 1;
        13'd1343: tone = `NM5 << 1;
        
        13'd1344: tone = `NM1 << 1;
        13'd1345: tone = `NM1 << 1;
        13'd1346: tone = `NM1 << 1;
        13'd1347: tone = `NM1 << 1;
        13'd1348: tone = `NM1 << 1;
        13'd1349: tone = `NM1 << 1;
        13'd1350: tone = `NM1 << 1;
        13'd1351: tone = `NM1 << 1;
        13'd1352: tone = `NM1 << 1;
        13'd1353: tone = `NM1 << 1;
        13'd1354: tone = `NM1 << 1;
        13'd1355: tone = `NM1 << 1;
        13'd1356: tone = `NM1 << 1;
        13'd1357: tone = `NM1 << 1;
        13'd1358: tone = `NM1 << 1;
        13'd1359: tone = `NM1 << 1;
        
        13'd1360: tone = `NM1 << 1;
        13'd1361: tone = `NM1 << 1;
        13'd1362: tone = `NM1 << 1;
        13'd1363: tone = `NM1 << 1;
        13'd1364: tone = `NM1 << 1;
        13'd1365: tone = `NM1 << 1;
        13'd1366: tone = `NM1 << 1;
        13'd1367: tone = `NM1 << 1;
        13'd1368: tone = `NM1 << 1;
        13'd1369: tone = `NM1 << 1;
        13'd1370: tone = `NM1 << 1;
        13'd1371: tone = `NM1 << 1;
        13'd1372: tone = `NM1 << 1;
        13'd1373: tone = `NM1 << 1;
        13'd1374: tone = `NM1 << 1;
        13'd1375: tone = `NM1 << 1;
        
        13'd1376: tone = `NM10;
        13'd1377: tone = `NM10;
        13'd1378: tone = `NM10;
        13'd1379: tone = `NM10;
        13'd1380: tone = `NM10;
        13'd1381: tone = `NM10;
        13'd1382: tone = `NM10;
        13'd1383: tone = `NM10;
        13'd1384: tone = `NM10;
        13'd1385: tone = `NM10;
        13'd1386: tone = `NM10;
        13'd1387: tone = `NM10;
        13'd1388: tone = `NM10;
        13'd1389: tone = `NM10;
        13'd1390: tone = `NM10;
        13'd1391: tone = `NM10;
        
        13'd1392: tone = `NM11;
        13'd1393: tone = `NM11;
        13'd1394: tone = `NM11;
        13'd1395: tone = `NM11;
        13'd1396: tone = `NM11;
        13'd1397: tone = `NM11;
        13'd1398: tone = `NM11;
        13'd1399: tone = `NM0;
        13'd1400: tone = `NM11;
        13'd1401: tone = `NM11;
        13'd1402: tone = `NM11;
        13'd1403: tone = `NM11;
        13'd1404: tone = `NM2 << 1;
        13'd1405: tone = `NM2 << 1;
        13'd1406: tone = `NM2 << 1;
        13'd1407: tone = `NM2 << 1;
        
        13'd1408: tone = `NM4 << 1;
        13'd1409: tone = `NM4 << 1;
        13'd1410: tone = `NM4 << 1;
        13'd1411: tone = `NM4 << 1;
        13'd1412: tone = `NM4 << 1;
        13'd1413: tone = `NM4 << 1;
        13'd1414: tone = `NM4 << 1;
        13'd1415: tone = `NM4 << 1;
        13'd1416: tone = `NM4 << 1;
        13'd1417: tone = `NM4 << 1;
        13'd1418: tone = `NM4 << 1;
        13'd1419: tone = `NM4 << 1;
        13'd1420: tone = `NM4 << 1;
        13'd1421: tone = `NM4 << 1;
        13'd1422: tone = `NM4 << 1;
        13'd1423: tone = `NM4 << 1;
        
        13'd1424: tone = `NM4 << 1;
        13'd1425: tone = `NM4 << 1;
        13'd1426: tone = `NM4 << 1;
        13'd1427: tone = `NM4 << 1;
        13'd1428: tone = `NM4 << 1;
        13'd1429: tone = `NM4 << 1;
        13'd1430: tone = `NM4 << 1;
        13'd1431: tone = `NM4 << 1;
        13'd1432: tone = `NM4 << 1;
        13'd1433: tone = `NM4 << 1;
        13'd1434: tone = `NM4 << 1;
        13'd1435: tone = `NM4 << 1;
        13'd1436: tone = `NM4 << 1;
        13'd1437: tone = `NM4 << 1;
        13'd1438: tone = `NM4 << 1;
        13'd1439: tone = `NM4 << 1;
        
        13'd1440: tone = `NM7 << 1;
        13'd1441: tone = `NM7 << 1;
        13'd1442: tone = `NM7 << 1;
        13'd1443: tone = `NM7 << 1;
        13'd1444: tone = `NM7 << 1;
        13'd1445: tone = `NM7 << 1;
        13'd1446: tone = `NM7 << 1;
        13'd1447: tone = `NM7 << 1;
        13'd1448: tone = `NM7 << 1;
        13'd1449: tone = `NM7 << 1;
        13'd1450: tone = `NM7 << 1;
        13'd1451: tone = `NM7 << 1;
        13'd1452: tone = `NM7 << 1;
        13'd1453: tone = `NM7 << 1;
        13'd1454: tone = `NM7 << 1;
        13'd1455: tone = `NM7 << 1;
        
        13'd1456: tone = `NM5 << 1;
        13'd1457: tone = `NM5 << 1;
        13'd1458: tone = `NM5 << 1;
        13'd1459: tone = `NM5 << 1;
        13'd1460: tone = `NM5 << 1;
        13'd1461: tone = `NM5 << 1;
        13'd1462: tone = `NM5 << 1;
        13'd1463: tone = `NM5 << 1;
        13'd1464: tone = `NM5;
        13'd1465: tone = `NM5;
        13'd1466: tone = `NM5;
        13'd1467: tone = `NM0;
        13'd1468: tone = `NM5;
        13'd1469: tone = `NM5;
        13'd1470: tone = `NM5;
        13'd1471: tone = `NM0;
        
        13'd1472: tone = `NM5;
        13'd1473: tone = `NM5;
        13'd1474: tone = `NM5;
        13'd1475: tone = `NM5;
        13'd1476: tone = `NM5;
        13'd1477: tone = `NM5;
        13'd1478: tone = `NM5;
        13'd1479: tone = `NM0;
        13'd1480: tone = `NM5;
        13'd1481: tone = `NM5;
        13'd1482: tone = `NM5;
        13'd1483: tone = `NM0;
        13'd1484: tone = `NM5;
        13'd1485: tone = `NM5;
        13'd1486: tone = `NM5;
        13'd1487: tone = `NM0;
        
        13'd1488: tone = `NM5;
        13'd1489: tone = `NM5;
        13'd1490: tone = `NM5;
        13'd1491: tone = `NM5;
        13'd1492: tone = `NM5;
        13'd1493: tone = `NM5;
        13'd1494: tone = `NM5;
        13'd1495: tone = `NM0;
        13'd1496: tone = `NM5;
        13'd1497: tone = `NM5;
        13'd1498: tone = `NM5;
        13'd1499: tone = `NM0;
        13'd1500: tone = `NM5;
        13'd1501: tone = `NM5;
        13'd1502: tone = `NM5;
        13'd1503: tone = `NM0;
        
        13'd1504: tone = `NM5;
        13'd1505: tone = `NM5;
        13'd1506: tone = `NM5;
        13'd1507: tone = `NM5;
        13'd1508: tone = `NM5;
        13'd1509: tone = `NM5;
        13'd1510: tone = `NM5;
        13'd1511: tone = `NM0;
        13'd1512: tone = `NM5;
        13'd1513: tone = `NM5;
        13'd1514: tone = `NM5;
        13'd1515: tone = `NM5;
        13'd1516: tone = `NM5;
        13'd1517: tone = `NM5;
        13'd1518: tone = `NM5;
        13'd1519: tone = `NM5;
		default : tone = `NM0;



	endcase
end

endmodule