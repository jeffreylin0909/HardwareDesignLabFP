//
//
//
//

`define NM1 32'd261 //C_freq
`define NM2 32'd277 //C#_freq
`define NM3 32'd294 //D_freq
`define NM4 32'd311 //Eb_freq
`define NM5 32'd330 //E_freq
`define NM6 32'd349 //F_freq
`define NM7 32'd370 //F#_freq
`define NM8 32'd392 //G_freq
`define NM9 32'd415 //G#_freq
`define NM10 32'd440 //A_freq
`define NM11 32'd466 //Bb_freq
`define NM12 32'd494 //B_freq
`define NM0 32'd20000 //slience (over freq.)

module MusicBoss (
	input [12:0] ibeatNum,	
	output reg [31:0] tone
);
//each block = 1 beat or quarter note
always @(*) begin
	case (ibeatNum)		// 1/16 beat 
		13'd0 : tone = `NM11 << 1;	
		13'd1 : tone = `NM11 << 1;
		13'd2 : tone = `NM11 << 1;
		13'd3 : tone = `NM11 << 1;
		13'd4 : tone = `NM11 << 1;	
		13'd5 : tone = `NM11 << 1;
		13'd6 : tone = `NM11 << 1;
		13'd7 : tone = `NM11 << 1;
		13'd8 : tone = `NM8 << 1;	
		13'd9 : tone = `NM8 << 1;
		13'd10 : tone = `NM8 << 1;
		13'd11 : tone = `NM8 << 1;
		13'd12 : tone = `NM8 << 1;	
		13'd13 : tone = `NM8 << 1;
		13'd14 : tone = `NM8 << 1;
		13'd15 : tone = `NM8 << 1;
		
		13'd16 : tone = `NM2 << 2;
		13'd17 : tone = `NM2 << 2;
		13'd18 : tone = `NM2 << 2;
		13'd19 : tone = `NM2 << 2;
		13'd20 : tone = `NM2 << 2;
		13'd21 : tone = `NM2 << 2;
		13'd22 : tone = `NM2 << 2;
		13'd23 : tone = `NM2 << 2;
		13'd24 : tone = `NM2 << 2;
		13'd25 : tone = `NM2 << 2;
		13'd26 : tone = `NM2 << 2;
		13'd27 : tone = `NM2 << 2;
		13'd28 : tone = `NM2 << 2;
		13'd29 : tone = `NM2 << 2;
		13'd30 : tone = `NM2 << 2;
		13'd31 : tone = `NM2 << 2;
		
		13'd32 : tone = `NM2 << 2;
		13'd33 : tone = `NM2 << 2;
		13'd34 : tone = `NM2 << 2;
		13'd35 : tone = `NM2 << 2;
		13'd36 : tone = `NM2 << 2;
		13'd37 : tone = `NM2 << 2;
		13'd38 : tone = `NM2 << 2;
		13'd39 : tone = `NM2 << 2;
		13'd40 : tone = `NM2 << 2;
		13'd41 : tone = `NM2 << 2;
		13'd42 : tone = `NM2 << 2;
		13'd43 : tone = `NM2 << 2;
		13'd44 : tone = `NM2 << 2;
		13'd45 : tone = `NM2 << 2;
		13'd46 : tone = `NM2 << 2;
		13'd47 : tone = `NM2 << 2;
		
		13'd48 : tone = `NM2 << 2;
		13'd49 : tone = `NM2 << 2;
		13'd50 : tone = `NM2 << 2;
		13'd51 : tone = `NM2 << 2;
		13'd52 : tone = `NM2 << 2;
		13'd53 : tone = `NM2 << 2;
		13'd54 : tone = `NM2 << 2;
		13'd55 : tone = `NM2 << 2;
		13'd56 : tone = `NM2 << 2;
		13'd57 : tone = `NM2 << 2;
		13'd58 : tone = `NM2 << 2;
		13'd59 : tone = `NM2 << 2;
		13'd60 : tone = `NM2 << 2;
		13'd61 : tone = `NM2 << 2;
		13'd62 : tone = `NM2 << 2;
		13'd63 : tone = `NM2 << 2;
		
		13'd64 : tone = `NM2 << 2;
		13'd65 : tone = `NM2 << 2;
		13'd66 : tone = `NM2 << 2;
		13'd67 : tone = `NM2 << 2;
		13'd68 : tone = `NM2 << 2;
		13'd69 : tone = `NM2 << 2;
		13'd70 : tone = `NM2 << 2;
		13'd71 : tone = `NM2 << 2;
		13'd72 : tone = `NM0;
		13'd73 : tone = `NM0;
		13'd74 : tone = `NM0;
		13'd75 : tone = `NM0;
		13'd76 : tone = `NM0;
		13'd77 : tone = `NM0;
		13'd78 : tone = `NM0;
		13'd79 : tone = `NM0;
		
		13'd80 : tone = `NM11 << 1;
		13'd81 : tone = `NM11 << 1;
		13'd82 : tone = `NM11 << 1;
		13'd83 : tone = `NM11 << 1;
		13'd84 : tone = `NM11 << 1;
		13'd85 : tone = `NM11 << 1;
		13'd86 : tone = `NM11 << 1;
		13'd87 : tone = `NM11 << 1;
		13'd88 : tone = `NM8 << 1;
		13'd89 : tone = `NM8 << 1;
		13'd90 : tone = `NM8 << 1;
		13'd91 : tone = `NM8 << 1;
		13'd92 : tone = `NM8 << 1;
		13'd93 : tone = `NM8 << 1;
		13'd94 : tone = `NM8 << 1;
		13'd95 : tone = `NM8 << 1;
		
		13'd96: tone = `NM2 << 2;
        13'd97: tone = `NM2 << 2;
        13'd98: tone = `NM2 << 2;
        13'd99: tone = `NM2 << 2;
        13'd100: tone = `NM2 << 2;
        13'd101: tone = `NM2 << 2;
        13'd102: tone = `NM2 << 2;
        13'd103: tone = `NM2 << 2;
        13'd104: tone = `NM2 << 2;
        13'd105: tone = `NM2 << 2;
        13'd106: tone = `NM2 << 2;
        13'd107: tone = `NM2 << 2;
        13'd108: tone = `NM0 << 2;
        13'd109: tone = `NM0 << 2;
        13'd110: tone = `NM0 << 2;
        13'd111: tone = `NM0 << 2;
        
        13'd112: tone = `NM2 << 2;
        13'd113: tone = `NM2 << 2;
        13'd114: tone = `NM2 << 2;
        13'd115: tone = `NM2 << 2;
        13'd116: tone = `NM2 << 2;
        13'd117: tone = `NM2 << 2;
        13'd118: tone = `NM2 << 2;
        13'd119: tone = `NM2 << 2;
        13'd120: tone = `NM2 << 2;
        13'd121: tone = `NM2 << 2;
        13'd122: tone = `NM2 << 2;
        13'd123: tone = `NM2 << 2;
        13'd124: tone = `NM0 << 2;
        13'd125: tone = `NM0 << 2;
        13'd126: tone = `NM0 << 2;
        13'd127: tone = `NM0 << 2;
		//1
		13'd128: tone = `NM3 << 2;
        13'd129: tone = `NM3 << 2;
        13'd130: tone = `NM3 << 2;
        13'd131: tone = `NM3 << 2;
        13'd132: tone = `NM3 << 2;
        13'd133: tone = `NM3 << 2;
        13'd134: tone = `NM3 << 2;
        13'd135: tone = `NM3 << 2;
        13'd136: tone = `NM3 << 2;
        13'd137: tone = `NM3 << 2;
        13'd138: tone = `NM3 << 2;
        13'd139: tone = `NM3 << 2;
        13'd140: tone = `NM3 << 2;
        13'd141: tone = `NM3 << 2;
        13'd142: tone = `NM3 << 2;
        13'd143: tone = `NM3 << 2;
        //2
        13'd144: tone = `NM3 << 2;
        13'd145: tone = `NM3 << 2;
        13'd146: tone = `NM3 << 2;
        13'd147: tone = `NM3 << 2;
        13'd148: tone = `NM3 << 2;
        13'd149: tone = `NM3 << 2;
        13'd150: tone = `NM3 << 2;
        13'd151: tone = `NM3 << 2;
        13'd152: tone = `NM3 << 2;
        13'd153: tone = `NM3 << 2;
        13'd154: tone = `NM3 << 2;
        13'd155: tone = `NM3 << 2;
        13'd156: tone = `NM3 << 2;
        13'd157: tone = `NM3 << 2;
        13'd158: tone = `NM3 << 2;
        13'd159: tone = `NM3 << 2;
        //3
        13'd160: tone = `NM3 << 2;
        13'd161: tone = `NM3 << 2;
        13'd162: tone = `NM3 << 2;
        13'd163: tone = `NM3 << 2;
        13'd164: tone = `NM3 << 2;
        13'd165: tone = `NM3 << 2;
        13'd166: tone = `NM3 << 2;
        13'd167: tone = `NM3 << 2;
        13'd168: tone = `NM3 << 2;
        13'd169: tone = `NM3 << 2;
        13'd170: tone = `NM3 << 2;
        13'd171: tone = `NM3 << 2;
        13'd172: tone = `NM3 << 2;
        13'd173: tone = `NM3 << 2;
        13'd174: tone = `NM3 << 2;
        13'd175: tone = `NM3 << 2;
        //4
        13'd176: tone = `NM3 << 2;
        13'd177: tone = `NM3 << 2;
        13'd178: tone = `NM3 << 2;
        13'd179: tone = `NM3 << 2;
        13'd180: tone = `NM3 << 2;
        13'd181: tone = `NM3 << 2;
        13'd182: tone = `NM3 << 2;
        13'd183: tone = `NM3 << 2;
        13'd184: tone = `NM3 << 2;
        13'd185: tone = `NM3 << 2;
        13'd186: tone = `NM3 << 2;
        13'd187: tone = `NM3 << 2;
        13'd188: tone = `NM3 << 2;
        13'd189: tone = `NM3 << 2;
        13'd190: tone = `NM3 << 2;
        13'd191: tone = `NM3 << 2;
		//5
		13'd192: tone = `NM3 << 2;
        13'd193: tone = `NM3 << 2;
        13'd194: tone = `NM3 << 2;
        13'd195: tone = `NM3 << 2;
        13'd196: tone = `NM3 << 2;
        13'd197: tone = `NM3 << 2;
        13'd198: tone = `NM3 << 2;
        13'd199: tone = `NM3 << 2;
        13'd200: tone = `NM3 << 2;
        13'd201: tone = `NM3 << 2;
        13'd202: tone = `NM3 << 2;
        13'd203: tone = `NM3 << 2;
        13'd204: tone = `NM3 << 2;
        13'd205: tone = `NM3 << 2;
        13'd206: tone = `NM3 << 2;
        13'd207: tone = `NM3 << 2;
        //6
        13'd208: tone = `NM3 << 2;
        13'd209: tone = `NM3 << 2;
        13'd210: tone = `NM3 << 2;
        13'd211: tone = `NM3 << 2;
        13'd212: tone = `NM3 << 2;
        13'd213: tone = `NM3 << 2;
        13'd214: tone = `NM3 << 2;
        13'd215: tone = `NM3 << 2;
        13'd216: tone = `NM3 << 2;
        13'd217: tone = `NM3 << 2;
        13'd218: tone = `NM3 << 2;
        13'd219: tone = `NM3 << 2;
        13'd220: tone = `NM3 << 2;
        13'd221: tone = `NM3 << 2;
        13'd222: tone = `NM3 << 2;
        13'd223: tone = `NM3 << 2;
        //7
        13'd224: tone = `NM3 << 2;
        13'd225: tone = `NM3 << 2;
        13'd226: tone = `NM3 << 2;
        13'd227: tone = `NM3 << 2;
        13'd228: tone = `NM3 << 2;
        13'd229: tone = `NM3 << 2;
        13'd230: tone = `NM3 << 2;
        13'd231: tone = `NM3 << 2;
        13'd232: tone = `NM3 << 2;
        13'd233: tone = `NM3 << 2;
        13'd234: tone = `NM3 << 2;
        13'd235: tone = `NM3 << 2;
        13'd236: tone = `NM3 << 2;
        13'd237: tone = `NM3 << 2;
        13'd238: tone = `NM3 << 2;
        13'd239: tone = `NM3 << 2;
        //8
        13'd240: tone = `NM3 << 2;
        13'd241: tone = `NM3 << 2;
        13'd242: tone = `NM3 << 2;
        13'd243: tone = `NM3 << 2;
        13'd244: tone = `NM3 << 2;
        13'd245: tone = `NM3 << 2;
        13'd246: tone = `NM3 << 2;
        13'd247: tone = `NM3 << 2;
        13'd248: tone = `NM3 << 2;
        13'd249: tone = `NM3 << 2;
        13'd250: tone = `NM3 << 2;
        13'd251: tone = `NM3 << 2;
        13'd252: tone = `NM3 << 2;
        13'd253: tone = `NM3 << 2;
        13'd254: tone = `NM3 << 2;
        13'd255: tone = `NM3 << 2;

		13'd256: tone = `NM11 << 1;
        13'd257: tone = `NM11 << 1;
        13'd258: tone = `NM11 << 1;
        13'd259: tone = `NM11 << 1;
        13'd260: tone = `NM11 << 1;
        13'd261: tone = `NM11 << 1;
        13'd262: tone = `NM11 << 1;
        13'd263: tone = `NM11 << 1;
        13'd264: tone = `NM8 << 1;
        13'd265: tone = `NM8 << 1;
        13'd266: tone = `NM8 << 1;
        13'd267: tone = `NM8 << 1;
        13'd268: tone = `NM8 << 1;
        13'd269: tone = `NM8 << 1;
        13'd270: tone = `NM8 << 1;
        13'd271: tone = `NM8 << 1;
        
        13'd272: tone = `NM2 << 2;
        13'd273: tone = `NM2 << 2;
        13'd274: tone = `NM2 << 2;
        13'd275: tone = `NM2 << 2;
        13'd276: tone = `NM2 << 2;
        13'd277: tone = `NM2 << 2;
        13'd278: tone = `NM2 << 2;
        13'd279: tone = `NM2 << 2;
        13'd280: tone = `NM2 << 2;
        13'd281: tone = `NM2 << 2;
        13'd282: tone = `NM2 << 2;
        13'd283: tone = `NM2 << 2;
        13'd284: tone = `NM2 << 2;
        13'd285: tone = `NM2 << 2;
        13'd286: tone = `NM2 << 2;
        13'd287: tone = `NM2 << 2;
        13'd288: tone = `NM2 << 2;
        13'd289: tone = `NM2 << 2;
        13'd290: tone = `NM2 << 2;
        13'd291: tone = `NM2 << 2;
        13'd292: tone = `NM2 << 2;
        13'd293: tone = `NM2 << 2;
        13'd294: tone = `NM2 << 2;
        13'd295: tone = `NM2 << 2;
        13'd296: tone = `NM2 << 2;
        13'd297: tone = `NM2 << 2;
        13'd298: tone = `NM2 << 2;
        13'd299: tone = `NM2 << 2;
        13'd300: tone = `NM2 << 2;
        13'd301: tone = `NM2 << 2;
        13'd302: tone = `NM2 << 2;
        13'd303: tone = `NM2 << 2;
        13'd304: tone = `NM2 << 2;
        13'd305: tone = `NM2 << 2;
        13'd306: tone = `NM2 << 2;
        13'd307: tone = `NM2 << 2;
        13'd308: tone = `NM2 << 2;
        13'd309: tone = `NM2 << 2;
        13'd310: tone = `NM2 << 2;
        13'd311: tone = `NM2 << 2;
        13'd312: tone = `NM2 << 2;
        13'd313: tone = `NM2 << 2;
        13'd314: tone = `NM2 << 2;
        13'd315: tone = `NM2 << 2;
        13'd316: tone = `NM2 << 2;
        13'd317: tone = `NM2 << 2;
        13'd318: tone = `NM2 << 2;
        13'd319: tone = `NM2 << 2;
        13'd320: tone = `NM2 << 2;
        13'd321: tone = `NM2 << 2;
        13'd322: tone = `NM2 << 2;
        13'd323: tone = `NM2 << 2;
        13'd324: tone = `NM2 << 2;
        13'd325: tone = `NM2 << 2;
        13'd326: tone = `NM2 << 2;
        13'd327: tone = `NM2 << 2;
        
        13'd328: tone = `NM0;
        13'd329: tone = `NM0;
        13'd330: tone = `NM0;
        13'd331: tone = `NM0;
        13'd332: tone = `NM0;
        13'd333: tone = `NM0;
        13'd334: tone = `NM0;
        13'd335: tone = `NM0;
        
        13'd336: tone = `NM11 << 1;
        13'd337: tone = `NM11 << 1;
        13'd338: tone = `NM11 << 1;
        13'd339: tone = `NM11 << 1;
        13'd340: tone = `NM11 << 1;
        13'd341: tone = `NM11 << 1;
        13'd342: tone = `NM11 << 1;
        13'd343: tone = `NM11 << 1;
        13'd344: tone = `NM8 << 1;
        13'd345: tone = `NM8 << 1;
        13'd346: tone = `NM8 << 1;
        13'd347: tone = `NM8 << 1;
        13'd348: tone = `NM8 << 1;
        13'd349: tone = `NM8 << 1;
        13'd350: tone = `NM8 << 1;
        13'd351: tone = `NM8 << 1;
        
        13'd352: tone = `NM2 << 2;
        13'd353: tone = `NM2 << 2;
        13'd354: tone = `NM2 << 2;
        13'd355: tone = `NM2 << 2;
        13'd356: tone = `NM2 << 2;
        13'd357: tone = `NM2 << 2;
        13'd358: tone = `NM2 << 2;
        13'd359: tone = `NM2 << 2;
        13'd360: tone = `NM2 << 2;
        13'd361: tone = `NM2 << 2;
        13'd362: tone = `NM2 << 2;
        13'd363: tone = `NM2 << 2;
        13'd364: tone = `NM0;
        13'd365: tone = `NM0;
        13'd366: tone = `NM0;
        13'd367: tone = `NM0;
        
        13'd368: tone = `NM2 << 2;
        13'd369: tone = `NM2 << 2;
        13'd370: tone = `NM2 << 2;
        13'd371: tone = `NM2 << 2;
        13'd372: tone = `NM2 << 2;
        13'd373: tone = `NM2 << 2;
        13'd374: tone = `NM2 << 2;
        13'd375: tone = `NM2 << 2;
        13'd376: tone = `NM2 << 2;
        13'd377: tone = `NM2 << 2;
        13'd378: tone = `NM2 << 2;
        13'd379: tone = `NM2 << 2;
        13'd380: tone = `NM0;
        13'd381: tone = `NM0;
        13'd382: tone = `NM0;
        13'd383: tone = `NM0;
        
        13'd384: tone = `NM3 << 2;
        13'd385: tone = `NM3 << 2;
        13'd386: tone = `NM3 << 2;
        13'd387: tone = `NM3 << 2;
        13'd388: tone = `NM3 << 2;
        13'd389: tone = `NM3 << 2;
        13'd390: tone = `NM3 << 2;
        13'd391: tone = `NM3 << 2;
        13'd392: tone = `NM3 << 2;
        13'd393: tone = `NM3 << 2;
        13'd394: tone = `NM3 << 2;
        13'd395: tone = `NM3 << 2;
        13'd396: tone = `NM3 << 2;
        13'd397: tone = `NM3 << 2;
        13'd398: tone = `NM3 << 2;
        13'd399: tone = `NM3 << 2;
        13'd400: tone = `NM3 << 2;
        13'd401: tone = `NM3 << 2;
        13'd402: tone = `NM3 << 2;
        13'd403: tone = `NM3 << 2;
        13'd404: tone = `NM3 << 2;
        13'd405: tone = `NM3 << 2;
        13'd406: tone = `NM3 << 2;
        13'd407: tone = `NM3 << 2;
        13'd408: tone = `NM3 << 2;
        13'd409: tone = `NM3 << 2;
        13'd410: tone = `NM3 << 2;
        13'd411: tone = `NM3 << 2;
        13'd412: tone = `NM3 << 2;
        13'd413: tone = `NM3 << 2;
        13'd414: tone = `NM3 << 2;
        13'd415: tone = `NM3 << 2;
        13'd416: tone = `NM3 << 2;
        13'd417: tone = `NM3 << 2;
        13'd418: tone = `NM3 << 2;
        13'd419: tone = `NM3 << 2;
        13'd420: tone = `NM3 << 2;
        13'd421: tone = `NM3 << 2;
        13'd422: tone = `NM3 << 2;
        13'd423: tone = `NM3 << 2;
        13'd424: tone = `NM3 << 2;
        13'd425: tone = `NM3 << 2;
        13'd426: tone = `NM3 << 2;
        13'd427: tone = `NM3 << 2;
        13'd428: tone = `NM3 << 2;
        13'd429: tone = `NM3 << 2;
        13'd430: tone = `NM3 << 2;
        13'd431: tone = `NM3 << 2;
        13'd432: tone = `NM3 << 2;
        13'd433: tone = `NM3 << 2;
        13'd434: tone = `NM3 << 2;
        13'd435: tone = `NM3 << 2;
        13'd436: tone = `NM3 << 2;
        13'd437: tone = `NM3 << 2;
        13'd438: tone = `NM3 << 2;
        13'd439: tone = `NM3 << 2;
        13'd440: tone = `NM3 << 2;
        13'd441: tone = `NM3 << 2;
        13'd442: tone = `NM3 << 2;
        13'd443: tone = `NM3 << 2;
        13'd444: tone = `NM3 << 2;
        13'd445: tone = `NM3 << 2;
        13'd446: tone = `NM3 << 2;
        13'd447: tone = `NM3 << 2;
        13'd448: tone = `NM3 << 2;
        13'd449: tone = `NM3 << 2;
        13'd450: tone = `NM3 << 2;
        13'd451: tone = `NM3 << 2;
        13'd452: tone = `NM3 << 2;
        13'd453: tone = `NM3 << 2;
        13'd454: tone = `NM3 << 2;
        13'd455: tone = `NM3 << 2;
        13'd456: tone = `NM3 << 2;
        13'd457: tone = `NM3 << 2;
        13'd458: tone = `NM3 << 2;
        13'd459: tone = `NM3 << 2;
        13'd460: tone = `NM3 << 2;
        13'd461: tone = `NM3 << 2;
        13'd462: tone = `NM3 << 2;
        13'd463: tone = `NM3 << 2;
        13'd464: tone = `NM3 << 2;
        13'd465: tone = `NM3 << 2;
        13'd466: tone = `NM3 << 2;
        13'd467: tone = `NM3 << 2;
        13'd468: tone = `NM3 << 2;
        13'd469: tone = `NM3 << 2;
        13'd470: tone = `NM3 << 2;
        13'd471: tone = `NM3 << 2;
        13'd472: tone = `NM3 << 2;
        13'd473: tone = `NM3 << 2;
        13'd474: tone = `NM3 << 2;
        13'd475: tone = `NM3 << 2;
        13'd476: tone = `NM3 << 2;
        13'd477: tone = `NM3 << 2;
        13'd478: tone = `NM3 << 2;
        13'd479: tone = `NM3 << 2;
        13'd480: tone = `NM3 << 2;
        13'd481: tone = `NM3 << 2;
        13'd482: tone = `NM3 << 2;
        13'd483: tone = `NM3 << 2;
        13'd484: tone = `NM3 << 2;
        13'd485: tone = `NM3 << 2;
        13'd486: tone = `NM3 << 2;
        13'd487: tone = `NM3 << 2;
        13'd488: tone = `NM3 << 2;
        13'd489: tone = `NM3 << 2;
        13'd490: tone = `NM3 << 2;
        13'd491: tone = `NM3 << 2;
        13'd492: tone = `NM3 << 2;
        13'd493: tone = `NM3 << 2;
        13'd494: tone = `NM3 << 2;
        13'd495: tone = `NM3 << 2;
        13'd496: tone = `NM3 << 2;
        13'd497: tone = `NM3 << 2;
        13'd498: tone = `NM3 << 2;
        13'd499: tone = `NM3 << 2;
        13'd500: tone = `NM3 << 2;
        13'd501: tone = `NM3 << 2;
        13'd502: tone = `NM3 << 2;
        13'd503: tone = `NM3 << 2;
        13'd504: tone = `NM3 << 2;
        13'd505: tone = `NM3 << 2;
        13'd506: tone = `NM3 << 2;
        13'd507: tone = `NM3 << 2;
        13'd508: tone = `NM3 << 2;
        13'd509: tone = `NM3 << 2;
        13'd510: tone = `NM3 << 2;
        13'd511: tone = `NM3 << 2;

        
        13'd512: tone = `NM0;
        13'd513: tone = `NM0;
        13'd514: tone = `NM0;
        13'd515: tone = `NM0;
        13'd516: tone = `NM0;
        13'd517: tone = `NM0;
        13'd518: tone = `NM0;
        13'd519: tone = `NM0;
        13'd520: tone = `NM0;
        13'd521: tone = `NM0;
        13'd522: tone = `NM0;
        13'd523: tone = `NM0;
        13'd524: tone = `NM0;
        13'd525: tone = `NM0;
        13'd526: tone = `NM0;
        13'd527: tone = `NM0;
        13'd528: tone = `NM0;
        13'd529: tone = `NM0;
        13'd530: tone = `NM0;
        13'd531: tone = `NM0;
        13'd532: tone = `NM0;
        13'd533: tone = `NM0;
        13'd534: tone = `NM0;
        13'd535: tone = `NM0;
        13'd536: tone = `NM0;
        13'd537: tone = `NM0;
        13'd538: tone = `NM0;
        13'd539: tone = `NM0;
        13'd540: tone = `NM0;
        13'd541: tone = `NM0;
        13'd542: tone = `NM0;
        13'd543: tone = `NM0;
        
        13'd544: tone = `NM4 << 1;
        13'd545: tone = `NM4 << 1;
        13'd546: tone = `NM4 << 1;
        13'd547: tone = `NM4 << 1;
        13'd548: tone = `NM4 << 1;
        13'd549: tone = `NM4 << 1;
        13'd550: tone = `NM4 << 1;
        13'd551: tone = `NM4 << 1;
        13'd552: tone = `NM4 << 1;
        13'd553: tone = `NM4 << 1;
        13'd554: tone = `NM4 << 1;
        13'd555: tone = `NM4 << 1;
        13'd556: tone = `NM4 << 1;
        13'd557: tone = `NM4 << 1;
        13'd558: tone = `NM4 << 1;
        13'd559: tone = `NM4 << 1;
        
        13'd560: tone = `NM0;
        13'd561: tone = `NM0;
        13'd562: tone = `NM0;
        13'd563: tone = `NM0;
        13'd564: tone = `NM0;
        13'd565: tone = `NM0;
        13'd566: tone = `NM0;
        13'd567: tone = `NM0;
        13'd568: tone = `NM1 << 1;
        13'd569: tone = `NM1 << 1;
        13'd570: tone = `NM1 << 1;
        13'd571: tone = `NM1 << 1;
        13'd572: tone = `NM1 << 1;
        13'd573: tone = `NM1 << 1;
        13'd574: tone = `NM1 << 1;
        13'd575: tone = `NM0;
        
       13'd576: tone = `NM3 << 1;
        13'd577: tone = `NM3 << 1;
        13'd578: tone = `NM3 << 1;
        13'd579: tone = `NM3 << 1;
        13'd580: tone = `NM3 << 1;
        13'd581: tone = `NM3 << 1;
        13'd582: tone = `NM3 << 1;
        13'd583: tone = `NM3 << 1;
        13'd584: tone = `NM3 << 1;
        13'd585: tone = `NM3 << 1;
        13'd586: tone = `NM3 << 1;
        13'd587: tone = `NM3 << 1;
        13'd588: tone = `NM3 << 1;
        13'd589: tone = `NM3 << 1;
        13'd590: tone = `NM3 << 1;
        13'd591: tone = `NM3 << 1;
        
        13'd592: tone = `NM0;
        13'd593: tone = `NM0;
        13'd594: tone = `NM0;
        13'd595: tone = `NM0;
        13'd596: tone = `NM0;
        13'd597: tone = `NM0;
        13'd598: tone = `NM0;
        13'd599: tone = `NM0;
        13'd600: tone = `NM0;
        13'd601: tone = `NM0;
        13'd602: tone = `NM0;
        13'd603: tone = `NM0;
        13'd604: tone = `NM0;
        13'd605: tone = `NM0;
        13'd606: tone = `NM0;
        13'd607: tone = `NM0;
        
        13'd608: tone = `NM1 << 1;
        13'd609: tone = `NM1 << 1;
        13'd610: tone = `NM1 << 1;
        13'd611: tone = `NM1 << 1;
        13'd612: tone = `NM1 << 1;
        13'd613: tone = `NM1 << 1;
        13'd614: tone = `NM1 << 1;
        13'd615: tone = `NM1 << 1;
        13'd616: tone = `NM1 << 1;
        13'd617: tone = `NM1 << 1;
        13'd618: tone = `NM1 << 1;
        13'd619: tone = `NM1 << 1;
        13'd620: tone = `NM1 << 1;
        13'd621: tone = `NM1 << 1;
        13'd622: tone = `NM1 << 1;
        13'd623: tone = `NM1 << 1;
        
        13'd624: tone = `NM0;
        13'd625: tone = `NM0;
        13'd626: tone = `NM0;
        13'd627: tone = `NM0;
        13'd628: tone = `NM0;
        13'd629: tone = `NM0;
        13'd630: tone = `NM0;
        13'd631: tone = `NM0;
        13'd632: tone = `NM10;
        13'd633: tone = `NM10;
        13'd634: tone = `NM10;
        13'd635: tone = `NM10;
        13'd636: tone = `NM10;
        13'd637: tone = `NM10;
        13'd638: tone = `NM10;
        13'd639: tone = `NM10;
        
        13'd640: tone = `NM11;
        13'd641: tone = `NM11;
        13'd642: tone = `NM11;
        13'd643: tone = `NM11;
        13'd644: tone = `NM11;
        13'd645: tone = `NM11;
        13'd646: tone = `NM11;
        13'd647: tone = `NM11;
        13'd648: tone = `NM11;
        13'd649: tone = `NM11;
        13'd650: tone = `NM11;
        13'd651: tone = `NM11;
        13'd652: tone = `NM11;
        13'd653: tone = `NM11;
        13'd654: tone = `NM11;
        13'd655: tone = `NM11;
        
        13'd656: tone = `NM0;
        13'd657: tone = `NM0;
        13'd658: tone = `NM0;
        13'd659: tone = `NM0;
        13'd660: tone = `NM0;
        13'd661: tone = `NM0;
        13'd662: tone = `NM0;
        13'd663: tone = `NM0;
        13'd664: tone = `NM0;
        13'd665: tone = `NM0;
        13'd666: tone = `NM0;
        13'd667: tone = `NM0;
        13'd668: tone = `NM0;
        13'd669: tone = `NM0;
        13'd670: tone = `NM0;
        13'd671: tone = `NM0;
        
        13'd672: tone = `NM10;
        13'd673: tone = `NM10;
        13'd674: tone = `NM10;
        13'd675: tone = `NM10;
        13'd676: tone = `NM10;
        13'd677: tone = `NM10;
        13'd678: tone = `NM10;
        13'd679: tone = `NM10;
        13'd680: tone = `NM10;
        13'd681: tone = `NM10;
        13'd682: tone = `NM10;
        13'd683: tone = `NM10;
        13'd684: tone = `NM10;
        13'd685: tone = `NM10;
        13'd686: tone = `NM10;
        13'd687: tone = `NM10;
        
        13'd688: tone = `NM0;
        13'd689: tone = `NM0;
        13'd690: tone = `NM0;
        13'd691: tone = `NM0;
        13'd692: tone = `NM0;
        13'd693: tone = `NM0;
        13'd694: tone = `NM0;
        13'd695: tone = `NM0;
        13'd696: tone = `NM7;
        13'd697: tone = `NM7;
        13'd698: tone = `NM7;
        13'd699: tone = `NM7;
        13'd700: tone = `NM7;
        13'd701: tone = `NM7;
        13'd702: tone = `NM7;
        13'd703: tone = `NM7;
        
        13'd704: tone = `NM8;
        13'd705: tone = `NM8;
        13'd706: tone = `NM8;
        13'd707: tone = `NM8;
        13'd708: tone = `NM8;
        13'd709: tone = `NM8;
        13'd710: tone = `NM8;
        13'd711: tone = `NM8;
        13'd712: tone = `NM8;
        13'd713: tone = `NM8;
        13'd714: tone = `NM8;
        13'd715: tone = `NM8;
        13'd716: tone = `NM8;
        13'd717: tone = `NM8;
        13'd718: tone = `NM8;
        13'd719: tone = `NM8;
        
        13'd720: tone = `NM11;
        13'd721: tone = `NM11;
        13'd722: tone = `NM11;
        13'd723: tone = `NM11;
        13'd724: tone = `NM11;
        13'd725: tone = `NM11;
        13'd726: tone = `NM11;
        13'd727: tone = `NM11;
        13'd728: tone = `NM11;
        13'd729: tone = `NM11;
        13'd730: tone = `NM11;
        13'd731: tone = `NM11;
        13'd732: tone = `NM11;
        13'd733: tone = `NM11;
        13'd734: tone = `NM11;
        13'd735: tone = `NM11;
        
        13'd736: tone = `NM3 << 1;
        13'd737: tone = `NM3 << 1;
        13'd738: tone = `NM3 << 1;
        13'd739: tone = `NM3 << 1;
        13'd740: tone = `NM3 << 1;
        13'd741: tone = `NM3 << 1;
        13'd742: tone = `NM3 << 1;
        13'd743: tone = `NM3 << 1;
        13'd744: tone = `NM3 << 1;
        13'd745: tone = `NM3 << 1;
        13'd746: tone = `NM3 << 1;
        13'd747: tone = `NM3 << 1;
        13'd748: tone = `NM3 << 1;
        13'd749: tone = `NM3 << 1;
        13'd750: tone = `NM3 << 1;
        13'd751: tone = `NM3 << 1;
        
        13'd752: tone = `NM4 << 1;
        13'd753: tone = `NM4 << 1;
        13'd754: tone = `NM4 << 1;
        13'd755: tone = `NM4 << 1;
        13'd756: tone = `NM4 << 1;
        13'd757: tone = `NM4 << 1;
        13'd758: tone = `NM4 << 1;
        13'd759: tone = `NM4 << 1;
        13'd760: tone = `NM4 << 1;
        13'd761: tone = `NM4 << 1;
        13'd762: tone = `NM4 << 1;
        13'd763: tone = `NM4 << 1;
        13'd764: tone = `NM4 << 1;
        13'd765: tone = `NM4 << 1;
        13'd766: tone = `NM4 << 1;
        13'd767: tone = `NM4 << 1;
        
        13'd768: tone = `NM0;
        13'd769: tone = `NM0;
        13'd770: tone = `NM0;
        13'd771: tone = `NM0;
        13'd772: tone = `NM0;
        13'd773: tone = `NM0;
        13'd774: tone = `NM0;
        13'd775: tone = `NM0;
        13'd776: tone = `NM8 << 1;
        13'd777: tone = `NM8 << 1;
        13'd778: tone = `NM8 << 1;
        13'd779: tone = `NM8 << 1;
        13'd780: tone = `NM8 << 1;
        13'd781: tone = `NM8 << 1;
        13'd782: tone = `NM8 << 1;
        13'd783: tone = `NM0;
        
        13'd784: tone = `NM8 << 1;
        13'd785: tone = `NM8 << 1;
        13'd786: tone = `NM8 << 1;
        13'd787: tone = `NM8 << 1;
        13'd788: tone = `NM8 << 1;
        13'd789: tone = `NM8 << 1;
        13'd790: tone = `NM8 << 1;
        13'd791: tone = `NM0;
        13'd792: tone = `NM8 << 1;
        13'd793: tone = `NM8 << 1;
        13'd794: tone = `NM8 << 1;
        13'd795: tone = `NM8 << 1;
        13'd796: tone = `NM8 << 1;
        13'd797: tone = `NM8 << 1;
        13'd798: tone = `NM8 << 1;
        13'd799: tone = `NM0;
        
        13'd800: tone = `NM8 << 1;
        13'd801: tone = `NM8 << 1;
        13'd802: tone = `NM8 << 1;
        13'd803: tone = `NM8 << 1;
        13'd804: tone = `NM8 << 1;
        13'd805: tone = `NM8 << 1;
        13'd806: tone = `NM8 << 1;
        13'd807: tone = `NM8 << 1;
        13'd808: tone = `NM8 << 1;
        13'd809: tone = `NM8 << 1;
        13'd810: tone = `NM8 << 1;
        13'd811: tone = `NM8 << 1;
        13'd812: tone = `NM8 << 1;
        13'd813: tone = `NM8 << 1;
        13'd814: tone = `NM8 << 1;
        13'd815: tone = `NM0;
        
        13'd816: tone = `NM8 << 1;
        13'd817: tone = `NM8 << 1;
        13'd818: tone = `NM8 << 1;
        13'd819: tone = `NM8 << 1;
        13'd820: tone = `NM8 << 1;
        13'd821: tone = `NM8 << 1;
        13'd822: tone = `NM8 << 1;
        13'd823: tone = `NM0;
        13'd824: tone = `NM8 << 1;
        13'd825: tone = `NM8 << 1;
        13'd826: tone = `NM8 << 1;
        13'd827: tone = `NM8 << 1;
        13'd828: tone = `NM8 << 1;
        13'd829: tone = `NM8 << 1;
        13'd830: tone = `NM8 << 1;
        13'd831: tone = `NM8 << 1;
        
        13'd832: tone = `NM11 << 1;
        13'd833: tone = `NM11 << 1;
        13'd834: tone = `NM11 << 1;
        13'd835: tone = `NM11 << 1;
        13'd836: tone = `NM11 << 1;
        13'd837: tone = `NM11 << 1;
        13'd838: tone = `NM11 << 1;
        13'd839: tone = `NM11 << 1;
        13'd840: tone = `NM8 << 1;
        13'd841: tone = `NM8 << 1;
        13'd842: tone = `NM8 << 1;
        13'd843: tone = `NM8 << 1;
        13'd844: tone = `NM8 << 1;
        13'd845: tone = `NM8 << 1;
        13'd846: tone = `NM8 << 1;
        13'd847: tone = `NM8 << 1;
        
        13'd848: tone = `NM11 << 1;
        13'd849: tone = `NM11 << 1;
        13'd850: tone = `NM11 << 1;
        13'd851: tone = `NM11 << 1;
        13'd852: tone = `NM11 << 1;
        13'd853: tone = `NM11 << 1;
        13'd854: tone = `NM11 << 1;
        13'd855: tone = `NM11 << 1;
        13'd856: tone = `NM8 << 1;
        13'd857: tone = `NM8 << 1;
        13'd858: tone = `NM8 << 1;
        13'd859: tone = `NM8 << 1;
        13'd860: tone = `NM8 << 1;
        13'd861: tone = `NM8 << 1;
        13'd862: tone = `NM8 << 1;
        13'd863: tone = `NM8 << 1;
        
        13'd864: tone = `NM11 << 1;
        13'd865: tone = `NM11 << 1;
        13'd866: tone = `NM11 << 1;
        13'd867: tone = `NM11 << 1;
        13'd868: tone = `NM11 << 1;
        13'd869: tone = `NM11 << 1;
        13'd870: tone = `NM11 << 1;
        13'd871: tone = `NM11 << 1;
        13'd872: tone = `NM11 << 1;
        13'd873: tone = `NM11 << 1;
        13'd874: tone = `NM11 << 1;
        13'd875: tone = `NM11 << 1;
        13'd876: tone = `NM11 << 1;
        13'd877: tone = `NM11 << 1;
        13'd878: tone = `NM11 << 1;
        13'd879: tone = `NM11 << 1;
        
        13'd880: tone = `NM8 << 1;
        13'd881: tone = `NM8 << 1;
        13'd882: tone = `NM8 << 1;
        13'd883: tone = `NM8 << 1;
        13'd884: tone = `NM8 << 1;
        13'd885: tone = `NM8 << 1;
        13'd886: tone = `NM8 << 1;
        13'd887: tone = `NM8 << 1;
        13'd888: tone = `NM8 << 1;
        13'd889: tone = `NM8 << 1;
        13'd890: tone = `NM8 << 1;
        13'd891: tone = `NM8 << 1;
        13'd892: tone = `NM8 << 1;
        13'd893: tone = `NM8 << 1;
        13'd894: tone = `NM8 << 1;
        13'd895: tone = `NM8 << 1;
        
        13'd896: tone = `NM0;
        13'd897: tone = `NM0;
        13'd898: tone = `NM0;
        13'd899: tone = `NM0;
        13'd900: tone = `NM0;
        13'd901: tone = `NM0;
        13'd902: tone = `NM0;
        13'd903: tone = `NM0;
        13'd904: tone = `NM8 << 1;
        13'd905: tone = `NM8 << 1;
        13'd906: tone = `NM8 << 1;
        13'd907: tone = `NM8 << 1;
        13'd908: tone = `NM8 << 1;
        13'd909: tone = `NM8 << 1;
        13'd910: tone = `NM8 << 1;
        13'd911: tone = `NM8 << 1;
        
        13'd912: tone = `NM8 << 1;
        13'd913: tone = `NM8 << 1;
        13'd914: tone = `NM8 << 1;
        13'd915: tone = `NM8 << 1;
        13'd916: tone = `NM8 << 1;
        13'd917: tone = `NM8 << 1;
        13'd918: tone = `NM8 << 1;
        13'd919: tone = `NM0;
        13'd920: tone = `NM8 << 1;
        13'd921: tone = `NM8 << 1;
        13'd922: tone = `NM8 << 1;
        13'd923: tone = `NM8 << 1;
        13'd924: tone = `NM8 << 1;
        13'd925: tone = `NM8 << 1;
        13'd926: tone = `NM8 << 1;
        13'd927: tone = `NM0;
        
        13'd928: tone = `NM7 << 1;
        13'd929: tone = `NM7 << 1;
        13'd930: tone = `NM7 << 1;
        13'd931: tone = `NM7 << 1;
        13'd932: tone = `NM7 << 1;
        13'd933: tone = `NM7 << 1;
        13'd934: tone = `NM7 << 1;
        13'd935: tone = `NM7 << 1;
        13'd936: tone = `NM7 << 1;
        13'd937: tone = `NM7 << 1;
        13'd938: tone = `NM7 << 1;
        13'd939: tone = `NM7 << 1;
        13'd940: tone = `NM7 << 1;
        13'd941: tone = `NM7 << 1;
        13'd942: tone = `NM7 << 1;
        13'd943: tone = `NM7 << 1;
        
        13'd944: tone = `NM7 << 1;
        13'd945: tone = `NM7 << 1;
        13'd946: tone = `NM7 << 1;
        13'd947: tone = `NM7 << 1;
        13'd948: tone = `NM7 << 1;
        13'd949: tone = `NM7 << 1;
        13'd950: tone = `NM7 << 1;
        13'd951: tone = `NM0;
        13'd952: tone = `NM7 << 1;
        13'd953: tone = `NM7 << 1;
        13'd954: tone = `NM7 << 1;
        13'd955: tone = `NM7 << 1;
        13'd956: tone = `NM7 << 1;
        13'd957: tone = `NM7 << 1;
        13'd958: tone = `NM7 << 1;
        13'd959: tone = `NM0;
        
        13'd960: tone = `NM3 << 1;
        13'd961: tone = `NM3 << 1;
        13'd962: tone = `NM3 << 1;
        13'd963: tone = `NM3 << 1;
        13'd964: tone = `NM3 << 1;
        13'd965: tone = `NM3 << 1;
        13'd966: tone = `NM3 << 1;
        13'd967: tone = `NM0;
        13'd968: tone = `NM3 << 1;
        13'd969: tone = `NM3 << 1;
        13'd970: tone = `NM3 << 1;
        13'd971: tone = `NM3 << 1;
        13'd972: tone = `NM3 << 1;
        13'd973: tone = `NM3 << 1;
        13'd974: tone = `NM3 << 1;
        13'd975: tone = `NM3 << 1;
        
        13'd976: tone = `NM4 << 1;
        13'd977: tone = `NM4 << 1;
        13'd978: tone = `NM4 << 1;
        13'd979: tone = `NM4 << 1;
        13'd980: tone = `NM4 << 1;
        13'd981: tone = `NM4 << 1;
        13'd982: tone = `NM4 << 1;
        13'd983: tone = `NM0;
        13'd984: tone = `NM4 << 1;
        13'd985: tone = `NM4 << 1;
        13'd986: tone = `NM4 << 1;
        13'd987: tone = `NM4<< 1;
        13'd988: tone = `NM4 << 1;
        13'd989: tone = `NM4 << 1;
        13'd990: tone = `NM4 << 1;
        13'd991: tone = `NM4 << 1;
        
        13'd992: tone = `NM3 << 1;
        13'd993: tone = `NM3 << 1;
        13'd994: tone = `NM3 << 1;
        13'd995: tone = `NM3 << 1;
        13'd996: tone = `NM3 << 1;
        13'd997: tone = `NM3 << 1;
        13'd998: tone = `NM3 << 1;
        13'd999: tone = `NM3 << 1;
        13'd1000: tone = `NM2 << 1;
        13'd1001: tone = `NM2 << 1;
        13'd1002: tone = `NM2 << 1;
        13'd1003: tone = `NM2 << 1;
        13'd1004: tone = `NM2 << 1;
        13'd1005: tone = `NM2 << 1;
        13'd1006: tone = `NM2 << 1;
        13'd1007: tone = `NM2 << 1;
        
        13'd1008: tone = `NM3 << 1;
        13'd1009: tone = `NM3 << 1;
        13'd1010: tone = `NM3 << 1;
        13'd1011: tone = `NM3 << 1;
        13'd1012: tone = `NM3 << 1;
        13'd1013: tone = `NM3 << 1;
        13'd1014: tone = `NM3 << 1;
        13'd1015: tone = `NM3 << 1;
        13'd1016: tone = `NM3 << 1;
        13'd1017: tone = `NM3 << 1;
        13'd1018: tone = `NM3 << 1;
        13'd1019: tone = `NM3 << 1;
        13'd1020: tone = `NM3 << 1;
        13'd1021: tone = `NM3 << 1;
        13'd1022: tone = `NM3 << 1;
        13'd1023: tone = `NM3 << 1;
        
       13'd1024: tone = `NM0;
        13'd1025: tone = `NM0;
        13'd1026: tone = `NM0;
        13'd1027: tone = `NM0;
        13'd1028: tone = `NM0;
        13'd1029: tone = `NM0;
        13'd1030: tone = `NM0;
        13'd1031: tone = `NM0;
        13'd1032: tone = `NM0;
        13'd1033: tone = `NM0;
        13'd1034: tone = `NM0;
        13'd1035: tone = `NM0;
        13'd1036: tone = `NM0;
        13'd1037: tone = `NM0;
        13'd1038: tone = `NM0;
        13'd1039: tone = `NM0;
        
        13'd1040: tone = `NM3 << 1;
        13'd1041: tone = `NM3 << 1;
        13'd1042: tone = `NM3 << 1;
        13'd1043: tone = `NM3 << 1;
        13'd1044: tone = `NM3 << 1;
        13'd1045: tone = `NM3 << 1;
        13'd1046: tone = `NM3 << 1;
        13'd1047: tone = `NM3 << 1;
        13'd1048: tone = `NM8;
        13'd1049: tone = `NM8;
        13'd1050: tone = `NM8;
        13'd1051: tone = `NM8;
        13'd1052: tone = `NM8;
        13'd1053: tone = `NM8;
        13'd1054: tone = `NM8;
        13'd1055: tone = `NM8;
        
        13'd1056: tone = `NM3 << 1;
        13'd1057: tone = `NM3 << 1;
        13'd1058: tone = `NM3 << 1;
        13'd1059: tone = `NM3 << 1;
        13'd1060: tone = `NM3 << 1;
        13'd1061: tone = `NM3 << 1;
        13'd1062: tone = `NM3 << 1;
        13'd1063: tone = `NM3 << 1;
        13'd1064: tone = `NM3 << 1;
        13'd1065: tone = `NM3 << 1;
        13'd1066: tone = `NM3 << 1;
        13'd1067: tone = `NM3 << 1;
        13'd1068: tone = `NM0;
        13'd1069: tone = `NM0;
        13'd1070: tone = `NM0;
        13'd1071: tone = `NM0;
        
        13'd1072: tone = `NM3 << 1;
        13'd1073: tone = `NM3 << 1;
        13'd1074: tone = `NM3 << 1;
        13'd1075: tone = `NM3 << 1;
        13'd1076: tone = `NM3 << 1;
        13'd1077: tone = `NM3 << 1;
        13'd1078: tone = `NM3 << 1;
        13'd1079: tone = `NM3 << 1;
        13'd1080: tone = `NM3 << 1;
        13'd1081: tone = `NM3 << 1;
        13'd1082: tone = `NM3 << 1;
        13'd1083: tone = `NM3 << 1;
        13'd1084: tone = `NM0;
        13'd1085: tone = `NM0;
        13'd1086: tone = `NM0;
        13'd1087: tone = `NM0;
        
        13'd1088: tone = `NM4 << 1;
        13'd1089: tone = `NM4 << 1;
        13'd1090: tone = `NM4 << 1;
        13'd1091: tone = `NM4 << 1;
        13'd1092: tone = `NM4 << 1;
        13'd1093: tone = `NM4 << 1;
        13'd1094: tone = `NM4 << 1;
        13'd1095: tone = `NM4 << 1;
        13'd1096: tone = `NM4 << 1;
        13'd1097: tone = `NM4 << 1;
        13'd1098: tone = `NM4 << 1;
        13'd1099: tone = `NM4 << 1;
        13'd1100: tone = `NM4 << 1;
        13'd1101: tone = `NM4 << 1;
        13'd1102: tone = `NM4 << 1;
        13'd1103: tone = `NM4 << 1;
        
        13'd1104: tone = `NM6 << 1;
        13'd1105: tone = `NM6 << 1;
        13'd1106: tone = `NM6 << 1;
        13'd1107: tone = `NM6 << 1;
        13'd1108: tone = `NM6 << 1;
        13'd1109: tone = `NM6 << 1;
        13'd1110: tone = `NM6 << 1;
        13'd1111: tone = `NM6 << 1;
        13'd1112: tone = `NM6 << 1;
        13'd1113: tone = `NM6 << 1;
        13'd1114: tone = `NM6 << 1;
        13'd1115: tone = `NM6 << 1;
        13'd1116: tone = `NM6 << 1;
        13'd1117: tone = `NM6 << 1;
        13'd1118: tone = `NM6 << 1;
        13'd1119: tone = `NM6 << 1;
        
        13'd1120: tone = `NM4 << 1;
        13'd1121: tone = `NM4 << 1;
        13'd1122: tone = `NM4 << 1;
        13'd1123: tone = `NM4 << 1;
        13'd1124: tone = `NM4 << 1;
        13'd1125: tone = `NM4 << 1;
        13'd1126: tone = `NM4 << 1;
        13'd1127: tone = `NM4 << 1;
        13'd1128: tone = `NM4 << 1;
        13'd1129: tone = `NM4 << 1;
        13'd1130: tone = `NM4 << 1;
        13'd1131: tone = `NM4 << 1;
        13'd1132: tone = `NM4 << 1;
        13'd1133: tone = `NM4 << 1;
        13'd1134: tone = `NM4 << 1;
        13'd1135: tone = `NM4 << 1;
        
        13'd1136: tone = `NM3 << 1;
        13'd1137: tone = `NM3 << 1;
        13'd1138: tone = `NM3 << 1;
        13'd1139: tone = `NM3 << 1;
        13'd1140: tone = `NM3 << 1;
        13'd1141: tone = `NM3 << 1;
        13'd1142: tone = `NM3 << 1;
        13'd1143: tone = `NM0;
        13'd1144: tone = `NM3 << 1;
        13'd1145: tone = `NM3 << 1;
        13'd1146: tone = `NM3 << 1;
        13'd1147: tone = `NM3 << 1;
        13'd1148: tone = `NM3 << 1;
        13'd1149: tone = `NM3 << 1;
        13'd1150: tone = `NM3 << 1;
        13'd1151: tone = `NM3 << 1;
        
        13'd1152: tone = `NM3 << 1;
        13'd1153: tone = `NM3 << 1;
        13'd1154: tone = `NM3 << 1;
        13'd1155: tone = `NM3 << 1;
        13'd1156: tone = `NM3 << 1;
        13'd1157: tone = `NM3 << 1;
        13'd1158: tone = `NM3 << 1;
        13'd1159: tone = `NM3 << 1;
        13'd1160: tone = `NM3 << 1;
        13'd1161: tone = `NM3 << 1;
        13'd1162: tone = `NM3 << 1;
        13'd1163: tone = `NM3 << 1;
        13'd1164: tone = `NM3 << 1;
        13'd1165: tone = `NM3 << 1;
        13'd1166: tone = `NM3 << 1;
        13'd1167: tone = `NM3 << 1;
        
        13'd1168: tone = `NM0;
        13'd1169: tone = `NM0;
        13'd1170: tone = `NM0;
        13'd1171: tone = `NM0;
        13'd1172: tone = `NM0;
        13'd1173: tone = `NM0;
        13'd1174: tone = `NM0;
        13'd1175: tone = `NM0;
        13'd1176: tone = `NM0;
        13'd1177: tone = `NM0;
        13'd1178: tone = `NM0;
        13'd1179: tone = `NM0;
        13'd1180: tone = `NM0;
        13'd1181: tone = `NM0;
        13'd1182: tone = `NM0;
        13'd1183: tone = `NM0;
        
        13'd1184: tone = `NM8 << 1;
        13'd1185: tone = `NM8 << 1;
        13'd1186: tone = `NM8 << 1;
        13'd1187: tone = `NM8 << 1;
        13'd1188: tone = `NM8 << 1;
        13'd1189: tone = `NM8 << 1;
        13'd1190: tone = `NM8 << 1;
        13'd1191: tone = `NM8 << 1;
        13'd1192: tone = `NM8 << 1;
        13'd1193: tone = `NM8 << 1;
        13'd1194: tone = `NM8 << 1;
        13'd1195: tone = `NM8 << 1;
        13'd1196: tone = `NM8 << 1;
        13'd1197: tone = `NM8 << 1;
        13'd1198: tone = `NM8 << 1;
        13'd1199: tone = `NM8 << 1;
        
        13'd1200: tone = `NM8 << 1;
        13'd1201: tone = `NM8 << 1;
        13'd1202: tone = `NM8 << 1;
        13'd1203: tone = `NM8 << 1;
        13'd1204: tone = `NM8 << 1;
        13'd1205: tone = `NM8 << 1;
        13'd1206: tone = `NM8 << 1;
        13'd1207: tone = `NM8 << 1;
        13'd1208: tone = `NM8 << 1;
        13'd1209: tone = `NM8 << 1;
        13'd1210: tone = `NM8 << 1;
        13'd1211: tone = `NM8 << 1;
        13'd1212: tone = `NM8 << 1;
        13'd1213: tone = `NM8 << 1;
        13'd1214: tone = `NM8 << 1;
        13'd1215: tone = `NM8 << 1;
        
        13'd1216: tone = `NM7 << 1;
        13'd1217: tone = `NM7 << 1;
        13'd1218: tone = `NM7 << 1;
        13'd1219: tone = `NM7 << 1;
        13'd1220: tone = `NM7 << 1;
        13'd1221: tone = `NM7 << 1;
        13'd1222: tone = `NM7 << 1;
        13'd1223: tone = `NM7 << 1;
        13'd1224: tone = `NM7 << 1;
        13'd1225: tone = `NM7 << 1;
        13'd1226: tone = `NM7 << 1;
        13'd1227: tone = `NM7 << 1;
        13'd1228: tone = `NM7 << 1;
        13'd1229: tone = `NM7 << 1;
        13'd1230: tone = `NM7 << 1;
        13'd1231: tone = `NM7 << 1;
        
        13'd1232: tone = `NM7 << 1;
        13'd1233: tone = `NM7 << 1;
        13'd1234: tone = `NM7 << 1;
        13'd1235: tone = `NM7 << 1;
        13'd1236: tone = `NM7 << 1;
        13'd1237: tone = `NM7 << 1;
        13'd1238: tone = `NM7 << 1;
        13'd1239: tone = `NM7 << 1;
        13'd1240: tone = `NM7 << 1;
        13'd1241: tone = `NM7 << 1;
        13'd1242: tone = `NM7 << 1;
        13'd1243: tone = `NM7 << 1;
        13'd1244: tone = `NM7 << 1;
        13'd1245: tone = `NM7 << 1;
        13'd1246: tone = `NM7 << 1;
        13'd1247: tone = `NM7 << 1;
        
        13'd1248: tone = `NM3 << 1;
        13'd1249: tone = `NM3 << 1;
        13'd1250: tone = `NM3 << 1;
        13'd1251: tone = `NM3 << 1;
        13'd1252: tone = `NM3 << 1;
        13'd1253: tone = `NM3 << 1;
        13'd1254: tone = `NM3 << 1;
        13'd1255: tone = `NM3 << 1;
        13'd1256: tone = `NM3 << 1;
        13'd1257: tone = `NM3 << 1;
        13'd1258: tone = `NM3 << 1;
        13'd1259: tone = `NM3 << 1;
        13'd1260: tone = `NM3 << 1;
        13'd1261: tone = `NM3 << 1;
        13'd1262: tone = `NM3 << 1;
        13'd1263: tone = `NM3 << 1;
        
        13'd1264: tone = `NM3 << 1;
        13'd1265: tone = `NM3 << 1;
        13'd1266: tone = `NM3 << 1;
        13'd1267: tone = `NM3 << 1;
        13'd1268: tone = `NM3 << 1;
        13'd1269: tone = `NM3 << 1;
        13'd1270: tone = `NM3 << 1;
        13'd1271: tone = `NM3 << 1;
        13'd1272: tone = `NM3 << 1;
        13'd1273: tone = `NM3 << 1;
        13'd1274: tone = `NM3 << 1;
        13'd1275: tone = `NM3 << 1;
        13'd1276: tone = `NM3 << 1;
        13'd1277: tone = `NM3 << 1;
        13'd1278: tone = `NM3 << 1;
        13'd1279: tone = `NM3 << 1;
        
        13'd1280: tone = `NM0;
        13'd1281: tone = `NM0;
        13'd1282: tone = `NM0;
        13'd1283: tone = `NM0;
        13'd1284: tone = `NM0;
        13'd1285: tone = `NM0;
        13'd1286: tone = `NM0;
        13'd1287: tone = `NM0;
        13'd1288: tone = `NM8 << 1;
        13'd1289: tone = `NM8 << 1;
        13'd1290: tone = `NM8 << 1;
        13'd1291: tone = `NM8 << 1;
        13'd1292: tone = `NM8 << 1;
        13'd1293: tone = `NM8 << 1;
        13'd1294: tone = `NM8 << 1;
        13'd1295: tone = `NM0;
        
        13'd1296: tone = `NM8 << 1;
        13'd1297: tone = `NM8 << 1;
        13'd1298: tone = `NM8 << 1;
        13'd1299: tone = `NM8 << 1;
        13'd1300: tone = `NM8 << 1;
        13'd1301: tone = `NM8 << 1;
        13'd1302: tone = `NM8 << 1;
        13'd1303: tone = `NM0;
        13'd1304: tone = `NM8 << 1;
        13'd1305: tone = `NM8 << 1;
        13'd1306: tone = `NM8 << 1;
        13'd1307: tone = `NM8 << 1;
        13'd1308: tone = `NM8 << 1;
        13'd1309: tone = `NM8 << 1;
        13'd1310: tone = `NM8 << 1;
        13'd1311: tone = `NM0;
        
        13'd1312: tone = `NM8 << 1;
        13'd1313: tone = `NM8 << 1;
        13'd1314: tone = `NM8 << 1;
        13'd1315: tone = `NM8 << 1;
        13'd1316: tone = `NM8 << 1;
        13'd1317: tone = `NM8 << 1;
        13'd1318: tone = `NM8 << 1;
        13'd1319: tone = `NM8 << 1;
        13'd1320: tone = `NM8 << 1;
        13'd1321: tone = `NM8 << 1;
        13'd1322: tone = `NM8 << 1;
        13'd1323: tone = `NM8 << 1;
        13'd1324: tone = `NM8 << 1;
        13'd1325: tone = `NM8 << 1;
        13'd1326: tone = `NM8 << 1;
        13'd1327: tone = `NM0;
        
        13'd1328: tone = `NM8 << 1;
        13'd1329: tone = `NM8 << 1;
        13'd1330: tone = `NM8 << 1;
        13'd1331: tone = `NM8 << 1;
        13'd1332: tone = `NM8 << 1;
        13'd1333: tone = `NM8 << 1;
        13'd1334: tone = `NM8 << 1;
        13'd1335: tone = `NM0 << 1;
        13'd1336: tone = `NM8 << 1;
        13'd1337: tone = `NM8 << 1;
        13'd1338: tone = `NM8 << 1;
        13'd1339: tone = `NM8 << 1;
        13'd1340: tone = `NM8 << 1;
        13'd1341: tone = `NM8 << 1;
        13'd1342: tone = `NM8 << 1;
        13'd1343: tone = `NM0;
        
        13'd1344: tone = `NM11 << 1;
        13'd1345: tone = `NM11 << 1;
        13'd1346: tone = `NM11 << 1;
        13'd1347: tone = `NM11 << 1;
        13'd1348: tone = `NM11 << 1;
        13'd1349: tone = `NM11 << 1;
        13'd1350: tone = `NM11 << 1;
        13'd1351: tone = `NM11 << 1;
        13'd1352: tone = `NM8 << 1;
        13'd1353: tone = `NM8 << 1;
        13'd1354: tone = `NM8 << 1;
        13'd1355: tone = `NM8 << 1;
        13'd1356: tone = `NM8 << 1;
        13'd1357: tone = `NM8 << 1;
        13'd1358: tone = `NM8 << 1;
        13'd1359: tone = `NM8 << 1;
        
        13'd1360: tone = `NM11 << 1;
        13'd1361: tone = `NM11 << 1;
        13'd1362: tone = `NM11 << 1;
        13'd1363: tone = `NM11 << 1;
        13'd1364: tone = `NM11 << 1;
        13'd1365: tone = `NM11 << 1;
        13'd1366: tone = `NM11 << 1;
        13'd1367: tone = `NM11 << 1;
        13'd1368: tone = `NM8 << 1;
        13'd1369: tone = `NM8 << 1;
        13'd1370: tone = `NM8 << 1;
        13'd1371: tone = `NM8 << 1;
        13'd1372: tone = `NM8 << 1;
        13'd1373: tone = `NM8 << 1;
        13'd1374: tone = `NM8 << 1;
        13'd1375: tone = `NM8 << 1;
        
        13'd1376: tone = `NM11 << 1;
        13'd1377: tone = `NM11 << 1;
        13'd1378: tone = `NM11 << 1;
        13'd1379: tone = `NM11 << 1;
        13'd1380: tone = `NM11 << 1;
        13'd1381: tone = `NM11 << 1;
        13'd1382: tone = `NM11 << 1;
        13'd1383: tone = `NM11 << 1;
        13'd1384: tone = `NM11 << 1;
        13'd1385: tone = `NM11 << 1;
        13'd1386: tone = `NM11 << 1;
        13'd1387: tone = `NM11 << 1;
        13'd1388: tone = `NM11 << 1;
        13'd1389: tone = `NM11 << 1;
        13'd1390: tone = `NM11 << 1;
        13'd1391: tone = `NM11 << 1;
        
        13'd1392: tone = `NM8 << 1;
        13'd1393: tone = `NM8 << 1;
        13'd1394: tone = `NM8 << 1;
        13'd1395: tone = `NM8 << 1;
        13'd1396: tone = `NM8 << 1;
        13'd1397: tone = `NM8 << 1;
        13'd1398: tone = `NM8 << 1;
        13'd1399: tone = `NM8 << 1;
        13'd1400: tone = `NM8 << 1;
        13'd1401: tone = `NM8 << 1;
        13'd1402: tone = `NM8 << 1;
        13'd1403: tone = `NM8 << 1;
        13'd1404: tone = `NM8 << 1;
        13'd1405: tone = `NM8 << 1;
        13'd1406: tone = `NM8 << 1;
        13'd1407: tone = `NM8 << 1;
        
        13'd1408: tone = `NM0;
        13'd1409: tone = `NM0;
        13'd1410: tone = `NM0;
        13'd1411: tone = `NM0;
        13'd1412: tone = `NM0;
        13'd1413: tone = `NM0;
        13'd1414: tone = `NM0;
        13'd1415: tone = `NM0;
        13'd1416: tone = `NM8 << 1;
        13'd1417: tone = `NM8 << 1;
        13'd1418: tone = `NM8 << 1;
        13'd1419: tone = `NM8 << 1;
        13'd1420: tone = `NM8 << 1;
        13'd1421: tone = `NM8 << 1;
        13'd1422: tone = `NM8 << 1;
        13'd1423: tone = `NM0;
        
        13'd1424: tone = `NM8 << 1;
        13'd1425: tone = `NM8 << 1;
        13'd1426: tone = `NM8 << 1;
        13'd1427: tone = `NM8 << 1;
        13'd1428: tone = `NM8 << 1;
        13'd1429: tone = `NM8 << 1;
        13'd1430: tone = `NM8 << 1;
        13'd1431: tone = `NM0;
        13'd1432: tone = `NM8 << 1;
        13'd1433: tone = `NM8 << 1;
        13'd1434: tone = `NM8 << 1;
        13'd1435: tone = `NM8 << 1;
        13'd1436: tone = `NM8 << 1;
        13'd1437: tone = `NM8 << 1;
        13'd1438: tone = `NM8 << 1;
        13'd1439: tone = `NM8 << 1;
        
        13'd1440: tone = `NM7 << 1;
        13'd1441: tone = `NM7 << 1;
        13'd1442: tone = `NM7 << 1;
        13'd1443: tone = `NM7 << 1;
        13'd1444: tone = `NM7 << 1;
        13'd1445: tone = `NM7 << 1;
        13'd1446: tone = `NM7 << 1;
        13'd1447: tone = `NM7 << 1;
        13'd1448: tone = `NM7 << 1;
        13'd1449: tone = `NM7 << 1;
        13'd1450: tone = `NM7 << 1;
        13'd1451: tone = `NM7 << 1;
        13'd1452: tone = `NM7 << 1;
        13'd1453: tone = `NM7 << 1;
        13'd1454: tone = `NM7 << 1;
        13'd1455: tone = `NM0;
        
        13'd1456: tone = `NM7 << 1;
        13'd1457: tone = `NM7 << 1;
        13'd1458: tone = `NM7 << 1;
        13'd1459: tone = `NM7 << 1;
        13'd1460: tone = `NM7 << 1;
        13'd1461: tone = `NM7 << 1;
        13'd1462: tone = `NM7 << 1;
        13'd1463: tone = `NM7 << 1;
        13'd1464: tone = `NM7 << 1;
        13'd1465: tone = `NM7 << 1;
        13'd1466: tone = `NM7 << 1;
        13'd1467: tone = `NM7 << 1;
        13'd1468: tone = `NM7 << 1;
        13'd1469: tone = `NM7 << 1;
        13'd1470: tone = `NM7 << 1;
        13'd1471: tone = `NM7 << 1;
        
        13'd1472: tone = `NM3 << 1;
        13'd1473: tone = `NM3 << 1;
        13'd1474: tone = `NM3 << 1;
        13'd1475: tone = `NM3 << 1;
        13'd1476: tone = `NM3 << 1;
        13'd1477: tone = `NM3 << 1;
        13'd1478: tone = `NM3 << 1;
        13'd1479: tone = `NM3 << 1;
        13'd1480: tone = `NM3 << 1;
        13'd1481: tone = `NM3 << 1;
        13'd1482: tone = `NM3 << 1;
        13'd1483: tone = `NM3 << 1;
        13'd1484: tone = `NM3 << 1;
        13'd1485: tone = `NM3 << 1;
        13'd1486: tone = `NM3 << 1;
        13'd1487: tone = `NM3 << 1;
        
        13'd1488: tone = `NM4 << 1;
        13'd1489: tone = `NM4 << 1;
        13'd1490: tone = `NM4 << 1;
        13'd1491: tone = `NM4 << 1;
        13'd1492: tone = `NM4 << 1;
        13'd1493: tone = `NM4 << 1;
        13'd1494: tone = `NM4 << 1;
        13'd1495: tone = `NM4 << 1;
        13'd1496: tone = `NM4 << 1;
        13'd1497: tone = `NM4 << 1;
        13'd1498: tone = `NM4 << 1;
        13'd1499: tone = `NM4 << 1;
        13'd1500: tone = `NM4 << 1;
        13'd1501: tone = `NM4 << 1;
        13'd1502: tone = `NM4 << 1;
        13'd1503: tone = `NM4 << 1;
        
        13'd1504: tone = `NM4 << 1;
        13'd1505: tone = `NM4 << 1;
        13'd1506: tone =  `NM4 << 1;
        13'd1507: tone = `NM4 << 1;
        13'd1508: tone = `NM4 << 1;
        13'd1509: tone = `NM4 << 1;
        13'd1510: tone = `NM4 << 1;
        13'd1511: tone = `NM4 << 1;
        13'd1512: tone = `NM0;
        13'd1513: tone = `NM0;
        13'd1514: tone = `NM0;
        13'd1515: tone = `NM0;
        13'd1516: tone = `NM0;
        13'd1517: tone = `NM0;
        13'd1518: tone = `NM0;
        13'd1519: tone = `NM0;
        
        13'd1520: tone = `NM2<< 1;
        13'd1521: tone = `NM2<< 1;
        13'd1522: tone = `NM2<< 1;
        13'd1523: tone = `NM2<< 1;
        13'd1524: tone = `NM2<< 1;
        13'd1525: tone = `NM2<< 1;
        13'd1526: tone = `NM2<< 1;
        13'd1527: tone = `NM2<< 1;
        13'd1528: tone = `NM3<< 1;
        13'd1529: tone = `NM3<< 1;
        13'd1530: tone = `NM3<< 1;
        13'd1531: tone = `NM3<< 1;
        13'd1532: tone = `NM3<< 1;
        13'd1533: tone = `NM3<< 1;
        13'd1534: tone = `NM3<< 1;
        13'd1535: tone = `NM3<< 1;
        
        13'd1536: tone = `NM4<< 1;
        13'd1537: tone = `NM4<< 1;
        13'd1538: tone = `NM4<< 1;
        13'd1539: tone = `NM4<< 1;
        13'd1540: tone = `NM4<< 1;
        13'd1541: tone = `NM4<< 1;
        13'd1542: tone = `NM4<< 1;
        13'd1543: tone = `NM4<< 1;
        13'd1544: tone = `NM4<< 1;
        13'd1545: tone = `NM4<< 1;
        13'd1546: tone = `NM4<< 1;
        13'd1547: tone = `NM4<< 1;
        13'd1548: tone = `NM4<< 1;
        13'd1549: tone = `NM4<< 1;
        13'd1550: tone = `NM4<< 1;
        13'd1551: tone = `NM4<< 1;
        
        13'd1552: tone = `NM3<< 1;
        13'd1553: tone = `NM3<< 1;
        13'd1554: tone = `NM3<< 1;
        13'd1555: tone = `NM3<< 1;
        13'd1556: tone = `NM3<< 1;
        13'd1557: tone = `NM3<< 1;
        13'd1558: tone = `NM3<< 1;
        13'd1559: tone = `NM3<< 1;
        13'd1560: tone = `NM2<<1;
        13'd1561: tone = `NM2<<1;
        13'd1562: tone = `NM2<<1;
        13'd1563: tone = `NM2<<1;
        13'd1564: tone = `NM2<<1;
        13'd1565: tone = `NM2<<1;
        13'd1566: tone = `NM2<<1;
        13'd1567: tone = `NM2<<1;
        
        13'd1568: tone = `NM3<< 1;
        13'd1569: tone = `NM3<< 1;
        13'd1570: tone = `NM3<< 1;
        13'd1571: tone = `NM3<< 1;
        13'd1572: tone = `NM3<< 1;
        13'd1573: tone = `NM3<< 1;
        13'd1574: tone = `NM3<< 1;
        13'd1575: tone = `NM3<< 1;
        13'd1576: tone = `NM2<<1;
        13'd1577: tone = `NM2<<1;
        13'd1578: tone = `NM2<<1;
        13'd1579: tone = `NM2<<1;
        13'd1580: tone = `NM2<<1;
        13'd1581: tone = `NM2<<1;
        13'd1582: tone = `NM2<<1;
        13'd1583: tone = `NM2<<1;
        
        13'd1584: tone = `NM3<<1;
        13'd1585: tone = `NM3<<1;
        13'd1586: tone = `NM3<<1;
        13'd1587: tone = `NM3<<1;
        13'd1588: tone = `NM3<<1;
        13'd1589: tone = `NM3<<1;
        13'd1590: tone = `NM3<<1;
        13'd1591: tone = `NM3<<1;
        13'd1592: tone = `NM3<<1;
        13'd1593: tone = `NM3<<1;
        13'd1594: tone = `NM3<<1;
        13'd1595: tone = `NM3<<1;
        13'd1596: tone = `NM3<<1;
        13'd1597: tone = `NM3<<1;
        13'd1598: tone = `NM3<<1;
        13'd1599: tone = `NM3<<1;
        
        13'd1600: tone = `NM3<<1;
        13'd1601: tone = `NM3<<1;
        13'd1602: tone = `NM3<<1;
        13'd1603: tone = `NM3<<1;
        13'd1604: tone = `NM3<<1;
        13'd1605: tone = `NM3<<1;
        13'd1606: tone = `NM3<<1;
        13'd1607: tone = `NM3<<1;
        13'd1608: tone = `NM3<<1;
        13'd1609: tone = `NM3<<1;
        13'd1610: tone = `NM3<<1;
        13'd1611: tone = `NM3<<1;
        13'd1612: tone = `NM3<<1;
        13'd1613: tone = `NM3<<1;
        13'd1614: tone = `NM3<<1;
        13'd1615: tone = `NM3<<1;
        
        13'd1616: tone = `NM3<<1;
        13'd1617: tone = `NM3<<1;
        13'd1618: tone = `NM3<<1;
        13'd1619: tone = `NM3<<1;
        13'd1620: tone = `NM3<<1;
        13'd1621: tone = `NM3<<1;
        13'd1622: tone = `NM3<<1;
        13'd1623: tone = `NM3<<1;
        13'd1624: tone = `NM3<<1;
        13'd1625: tone = `NM3<<1;
        13'd1626: tone = `NM3<<1;
        13'd1627: tone = `NM3<<1;
        13'd1628: tone = `NM3<<1;
        13'd1629: tone = `NM3<<1;
        13'd1630: tone = `NM3<<1;
        13'd1631: tone = `NM3<<1;
                
        13'd1632: tone = `NM0;
        13'd1633: tone = `NM0;
        13'd1634: tone = `NM0;
        13'd1635: tone = `NM0;
        13'd1636: tone = `NM0;
        13'd1637: tone = `NM0;
        13'd1638: tone = `NM0;
        13'd1639: tone = `NM0;
        13'd1640: tone = `NM0;
        13'd1641: tone = `NM0;
        13'd1642: tone = `NM0;
        13'd1643: tone = `NM0;
        13'd1644: tone = `NM0;
        13'd1645: tone = `NM0;
        13'd1646: tone = `NM0;
        13'd1647: tone = `NM0;
        
        13'd1648: tone = `NM2 << 1;
        13'd1649: tone = `NM2 << 1;
        13'd1650: tone = `NM2 << 1;
        13'd1651: tone = `NM2 << 1;
        13'd1652: tone = `NM2 << 1;
        13'd1653: tone = `NM2 << 1;
        13'd1654: tone = `NM2 << 1;
        13'd1655: tone = `NM2 << 1;
        13'd1656: tone = `NM3 << 1;
        13'd1657: tone = `NM3 << 1;
        13'd1658: tone = `NM3 << 1;
        13'd1659: tone = `NM3 << 1;
        13'd1660: tone = `NM3 << 1;
        13'd1661: tone = `NM3 << 1;
        13'd1662: tone = `NM3 << 1;
        13'd1663: tone = `NM3 << 1;
        
        13'd1664: tone = `NM3<<1;
        13'd1665: tone = `NM3<<1;
        13'd1666: tone = `NM3<<1;
        13'd1667: tone = `NM3<<1;
        13'd1668: tone = `NM3<<1;
        13'd1669: tone = `NM3<<1;
        13'd1670: tone = `NM3<<1;
        13'd1671: tone = `NM3<<1;
        13'd1672: tone = `NM3<<1;
        13'd1673: tone = `NM3<<1;
        13'd1674: tone = `NM3<<1;
        13'd1675: tone = `NM3<<1;
        13'd1676: tone = `NM3<<1;
        13'd1677: tone = `NM3<<1;
        13'd1678: tone = `NM3<<1;
        13'd1679: tone = `NM3<<1;
        
        13'd1680: tone = `NM3<<1;
        13'd1681: tone = `NM3<<1;
        13'd1682: tone = `NM3<<1;
        13'd1683: tone = `NM3<<1;
        13'd1684: tone = `NM3<<1;
        13'd1685: tone = `NM3<<1;
        13'd1686: tone = `NM3<<1;
        13'd1687: tone = `NM3<<1;
        13'd1688: tone = `NM3<<1;
        13'd1689: tone = `NM3<<1;
        13'd1690: tone = `NM3<<1;
        13'd1691: tone = `NM3<<1;
        13'd1692: tone = `NM3<<1;
        13'd1693: tone = `NM3<<1;
        13'd1694: tone = `NM3<<1;
        13'd1695: tone = `NM3<<1;
        
        13'd1696: tone = `NM3<<1;
        13'd1697: tone = `NM3<<1;
        13'd1698: tone = `NM3<<1;
        13'd1699: tone = `NM3<<1;
        13'd1700: tone = `NM3<<1;
        13'd1701: tone = `NM3<<1;
        13'd1702: tone = `NM3<<1;
        13'd1703: tone = `NM3<<1;
        13'd1704: tone = `NM3<<1;
        13'd1705: tone = `NM3<<1;
        13'd1706: tone = `NM3<<1;
        13'd1707: tone = `NM3<<1;
        13'd1708: tone = `NM3<<1;
        13'd1709: tone = `NM3<<1;
        13'd1710: tone = `NM3<<1;
        13'd1711: tone = `NM3<<1;
        
        13'd1712: tone = `NM3<<1;
        13'd1713: tone = `NM3<<1;
        13'd1714: tone = `NM3<<1;
        13'd1715: tone = `NM3<<1;
        13'd1716: tone = `NM3<<1;
        13'd1717: tone = `NM3<<1;
        13'd1718: tone = `NM3<<1;
        13'd1719: tone = `NM3<<1;
        13'd1720: tone = `NM3<<1;
        13'd1721: tone = `NM3<<1;
        13'd1722: tone = `NM3<<1;
        13'd1723: tone = `NM3<<1;
        13'd1724: tone = `NM3<<1;
        13'd1725: tone = `NM3<<1;
        13'd1726: tone = `NM3<<1;
        13'd1727: tone = `NM3<<1;
        
        13'd1728: tone = `NM3<<1;
        13'd1729: tone = `NM3<<1;
        13'd1730: tone = `NM3<<1;
        13'd1731: tone = `NM3<<1;
        13'd1732: tone = `NM3<<1;
        13'd1733: tone = `NM3<<1;
        13'd1734: tone = `NM3<<1;
        13'd1735: tone = `NM3<<1;
        13'd1736: tone = `NM3<<1;
        13'd1737: tone = `NM3<<1;
        13'd1738: tone = `NM3<<1;
        13'd1739: tone = `NM3<<1;
        13'd1740: tone = `NM3<<1;
        13'd1741: tone = `NM3<<1;
        13'd1742: tone = `NM3<<1;
        13'd1743: tone = `NM3<<1;
        
        13'd1744: tone = `NM3<<1;
        13'd1745: tone = `NM3<<1;
        13'd1746: tone = `NM3<<1;
        13'd1747: tone = `NM3<<1;
        13'd1748: tone = `NM3<<1;
        13'd1749: tone = `NM3<<1;
        13'd1750: tone = `NM3<<1;
        13'd1751: tone = `NM3<<1;
        13'd1752: tone = `NM3<<1;
        13'd1753: tone = `NM3<<1;
        13'd1754: tone = `NM3<<1;
        13'd1755: tone = `NM3<<1;
        13'd1756: tone = `NM3<<1;
        13'd1757: tone = `NM3<<1;
        13'd1758: tone = `NM3<<1;
        13'd1759: tone = `NM3<<1;
        
        13'd1760: tone = `NM0;
        13'd1761: tone = `NM0;
        13'd1762: tone = `NM0;
        13'd1763: tone = `NM0;
        13'd1764: tone = `NM0;
        13'd1765: tone = `NM0;
        13'd1766: tone = `NM0;
        13'd1767: tone = `NM0;
        13'd1768: tone = `NM0;
        13'd1769: tone = `NM0;
        13'd1770: tone = `NM0;
        13'd1771: tone = `NM0;
        13'd1772: tone = `NM0;
        13'd1773: tone = `NM0;
        13'd1774: tone = `NM0;
        13'd1775: tone = `NM0;
        
        13'd1776: tone = `NM2 << 1;
        13'd1777: tone = `NM2 << 1;
        13'd1778: tone = `NM2 << 1;
        13'd1779: tone = `NM2 << 1;
        13'd1780: tone = `NM2 << 1;
        13'd1781: tone = `NM2 << 1;
        13'd1782: tone = `NM2 << 1;
        13'd1783: tone = `NM2 << 1;
        13'd1784: tone = `NM3 << 1;
        13'd1785: tone = `NM3 << 1;
        13'd1786: tone = `NM3 << 1;
        13'd1787: tone = `NM3 << 1;
        13'd1788: tone = `NM3 << 1;
        13'd1789: tone = `NM3 << 1;
        13'd1790: tone = `NM3 << 1;
        13'd1791: tone = `NM3 << 1;
        
        13'd1792: tone = `NM4<<1;
        13'd1793: tone = `NM4<<1;
        13'd1794: tone = `NM4<<1;
        13'd1795: tone = `NM4<<1;
        13'd1796: tone = `NM4<<1;
        13'd1797: tone = `NM4<<1;
        13'd1798: tone = `NM4<<1;
        13'd1799: tone = `NM4<<1;
        13'd1800: tone = `NM4<<1;
        13'd1801: tone = `NM4<<1;
        13'd1802: tone = `NM4<<1;
        13'd1803: tone = `NM4<<1;
        13'd1804: tone = `NM4<<1;
        13'd1805: tone = `NM4<<1;
        13'd1806: tone = `NM4<<1;
        13'd1807: tone = `NM4<<1;
        
        13'd1808: tone = `NM3 << 1;
        13'd1809: tone = `NM3 << 1;
        13'd1810: tone = `NM3 << 1;
        13'd1811: tone = `NM3 << 1;
        13'd1812: tone = `NM3 << 1;
        13'd1813: tone = `NM3 << 1;
        13'd1814: tone = `NM3 << 1;
        13'd1815: tone = `NM3 << 1;
        13'd1816: tone = `NM2 << 1;
        13'd1817: tone = `NM2 << 1;
        13'd1818: tone = `NM2 << 1;
        13'd1819: tone = `NM2 << 1;
        13'd1820: tone = `NM2 << 1;
        13'd1821: tone = `NM2 << 1;
        13'd1822: tone = `NM2 << 1;
        13'd1823: tone = `NM2 << 1;
        
        13'd1824: tone = `NM3 << 1;
        13'd1825: tone = `NM3 << 1;
        13'd1826: tone = `NM3 << 1;
        13'd1827: tone = `NM3 << 1;
        13'd1828: tone = `NM3 << 1;
        13'd1829: tone = `NM3 << 1;
        13'd1830: tone = `NM3 << 1;
        13'd1831: tone = `NM3 << 1;
        13'd1832: tone = `NM2 << 1;
        13'd1833: tone = `NM2 << 1;
        13'd1834: tone = `NM2 << 1;
        13'd1835: tone = `NM2 << 1;
        13'd1836: tone = `NM2 << 1;
        13'd1837: tone = `NM2 << 1;
        13'd1838: tone = `NM2 << 1;
        13'd1839: tone = `NM2 << 1;
        
        13'd1840: tone = `NM3<<1;
        13'd1841: tone = `NM3<<1;
        13'd1842: tone = `NM3<<1;
        13'd1843: tone = `NM3<<1;
        13'd1844: tone = `NM3<<1;
        13'd1845: tone = `NM3<<1;
        13'd1846: tone = `NM3<<1;
        13'd1847: tone = `NM3<<1;
        13'd1848: tone = `NM3<<1;
        13'd1849: tone = `NM3<<1;
        13'd1850: tone = `NM3<<1;
        13'd1851: tone = `NM3<<1;
        13'd1852: tone = `NM3<<1;
        13'd1853: tone = `NM3<<1;
        13'd1854: tone = `NM3<<1;
        13'd1855: tone = `NM3<<1;
        
        13'd1856: tone = `NM3<<1;
        13'd1857: tone = `NM3<<1;
        13'd1858: tone = `NM3<<1;
        13'd1859: tone = `NM3<<1;
        13'd1860: tone = `NM3<<1;
        13'd1861: tone = `NM3<<1;
        13'd1862: tone = `NM3<<1;
        13'd1863: tone = `NM3<<1;
        13'd1864: tone = `NM3<<1;
        13'd1865: tone = `NM3<<1;
        13'd1866: tone = `NM3<<1;
        13'd1867: tone = `NM3<<1;
        13'd1868: tone = `NM3<<1;
        13'd1869: tone = `NM3<<1;
        13'd1870: tone = `NM3<<1;
        13'd1871: tone = `NM3<<1;
        
        13'd1872: tone = `NM3<<1;
        13'd1873: tone = `NM3<<1;
        13'd1874: tone = `NM3<<1;
        13'd1875: tone = `NM3<<1;
        13'd1876: tone = `NM3<<1;
        13'd1877: tone = `NM3<<1;
        13'd1878: tone = `NM3<<1;
        13'd1879: tone = `NM3<<1;
        13'd1880: tone = `NM3<<1;
        13'd1881: tone = `NM3<<1;
        13'd1882: tone = `NM3<<1;
        13'd1883: tone = `NM3<<1;
        13'd1884: tone = `NM3<<1;
        13'd1885: tone = `NM3<<1;
        13'd1886: tone = `NM3<<1;
        13'd1887: tone = `NM3<<1;
        
        13'd1888: tone = `NM0;
        13'd1889: tone = `NM0;
        13'd1890: tone = `NM0;
        13'd1891: tone = `NM0;
        13'd1892: tone = `NM0;
        13'd1893: tone = `NM0;
        13'd1894: tone = `NM0;
        13'd1895: tone = `NM0;
        13'd1896: tone = `NM0;
        13'd1897: tone = `NM0;
        13'd1898: tone = `NM0;
        13'd1899: tone = `NM0;
        13'd1900: tone = `NM0;
        13'd1901: tone = `NM0;
        13'd1902: tone = `NM0;
        13'd1903: tone = `NM0;
        
        13'd1904: tone = `NM7 << 1;
        13'd1905: tone = `NM7 << 1;
        13'd1906: tone = `NM7 << 1;
        13'd1907: tone = `NM7 << 1;
        13'd1908: tone = `NM7 << 1;
        13'd1909: tone = `NM7 << 1;
        13'd1910: tone = `NM7 << 1;
        13'd1911: tone = `NM7 << 1;
        13'd1912: tone = `NM8 << 1;
        13'd1913: tone = `NM8 << 1;
        13'd1914: tone = `NM8 << 1;
        13'd1915: tone = `NM8 << 1;
        13'd1916: tone = `NM8 << 1;
        13'd1917: tone = `NM8 << 1;
        13'd1918: tone = `NM8 << 1;
        13'd1919: tone = `NM8 << 1;
        
        13'd1920: tone = `NM8 << 1;
        13'd1921: tone = `NM8 << 1;
        13'd1922: tone = `NM8 << 1;
        13'd1923: tone = `NM8 << 1;
        13'd1924: tone = `NM8 << 1;
        13'd1925: tone = `NM8 << 1;
        13'd1926: tone = `NM8 << 1;
        13'd1927: tone = `NM8 << 1;
        13'd1928: tone = `NM8 << 1;
        13'd1929: tone = `NM8 << 1;
        13'd1930: tone = `NM8 << 1;
        13'd1931: tone = `NM8 << 1;
        13'd1932: tone = `NM8 << 1;
        13'd1933: tone = `NM8 << 1;
        13'd1934: tone = `NM8 << 1;
        13'd1935: tone = `NM8 << 1;
        
        13'd1936: tone = `NM8 << 1;
        13'd1937: tone = `NM8 << 1;
        13'd1938: tone = `NM8 << 1;
        13'd1939: tone = `NM8 << 1;
        13'd1940: tone = `NM8 << 1;
        13'd1941: tone = `NM8 << 1;
        13'd1942: tone = `NM8 << 1;
        13'd1943: tone = `NM8 << 1;
        13'd1944: tone = `NM8 << 1;
        13'd1945: tone = `NM8 << 1;
        13'd1946: tone = `NM8 << 1;
        13'd1947: tone = `NM8 << 1;
        13'd1948: tone = `NM8 << 1;
        13'd1949: tone = `NM8 << 1;
        13'd1950: tone = `NM8 << 1;
        13'd1951: tone = `NM8 << 1;
        
        13'd1952: tone = `NM8 << 1;
        13'd1953: tone = `NM8 << 1;
        13'd1954: tone = `NM8 << 1;
        13'd1955: tone = `NM8 << 1;
        13'd1956: tone = `NM8 << 1;
        13'd1957: tone = `NM8 << 1;
        13'd1958: tone = `NM8 << 1;
        13'd1959: tone = `NM8 << 1;
        13'd1960: tone = `NM8 << 1;
        13'd1961: tone = `NM8 << 1;
        13'd1962: tone = `NM8 << 1;
        13'd1963: tone = `NM8 << 1;
        13'd1964: tone = `NM8 << 1;
        13'd1965: tone = `NM8 << 1;
        13'd1966: tone = `NM8 << 1;
        13'd1967: tone = `NM8 << 1;
        
        13'd1968: tone = `NM8 << 1;
        13'd1969: tone = `NM8 << 1;
        13'd1970: tone = `NM8 << 1;
        13'd1971: tone = `NM8 << 1;
        13'd1972: tone = `NM8 << 1;
        13'd1973: tone = `NM8 << 1;
        13'd1974: tone = `NM8 << 1;
        13'd1975: tone = `NM8 << 1;
        13'd1976: tone = `NM8 << 1;
        13'd1977: tone = `NM8 << 1;
        13'd1978: tone = `NM8 << 1;
        13'd1979: tone = `NM8 << 1;
        13'd1980: tone = `NM8 << 1;
        13'd1981: tone = `NM8 << 1;
        13'd1982: tone = `NM8 << 1;
        13'd1983: tone = `NM8 << 1;
        
        13'd1984: tone = `NM0;
        13'd1985: tone = `NM0;
        13'd1986: tone = `NM0;
        13'd1987: tone = `NM0;
        13'd1988: tone = `NM0;
        13'd1989: tone = `NM0;
        13'd1990: tone = `NM0;
        13'd1991: tone = `NM0;
        13'd1992: tone = `NM0;
        13'd1993: tone = `NM0;
        13'd1994: tone = `NM0;
        13'd1995: tone = `NM0;
        13'd1996: tone = `NM0;
        13'd1997: tone = `NM0;
        13'd1998: tone = `NM0;
        13'd1999: tone = `NM0;
        
        13'd2000: tone = `NM0;
        13'd2001: tone = `NM0;
        13'd2002: tone = `NM0;
        13'd2003: tone = `NM0;
        13'd2004: tone = `NM0;
        13'd2005: tone = `NM0;
        13'd2006: tone = `NM0;
        13'd2007: tone = `NM0;
        13'd2008: tone = `NM8 << 1;
        13'd2009: tone = `NM8 << 1;
        13'd2010: tone = `NM8 << 1;
        13'd2011: tone = `NM8 << 1;
        13'd2012: tone = `NM8 << 1;
        13'd2013: tone = `NM8 << 1;
        13'd2014: tone = `NM8 << 1;
        13'd2015: tone = `NM8 << 1;
        
        13'd2016: tone = `NM11 <<1;
        13'd2017: tone = `NM11 <<1;
        13'd2018: tone = `NM11 <<1;
        13'd2019: tone = `NM11 <<1;
        13'd2020: tone = `NM11 <<1;
        13'd2021: tone = `NM11 <<1;
        13'd2022: tone = `NM11 <<1;
        13'd2023: tone = `NM0;
        13'd2024: tone = `NM11 <<1;
        13'd2025: tone = `NM11 <<1;
        13'd2026: tone = `NM11 <<1;
        13'd2027: tone = `NM11 <<1;
        13'd2028: tone = `NM11 <<1;
        13'd2029: tone = `NM11 <<1;
        13'd2030: tone = `NM11 <<1;
        13'd2031: tone = `NM0;
        
        13'd2032: tone = `NM8 << 1;
        13'd2033: tone = `NM8 << 1;
        13'd2034: tone = `NM8 << 1;
        13'd2035: tone = `NM8 << 1;
        13'd2036: tone = `NM8 << 1;
        13'd2037: tone = `NM8 << 1;
        13'd2038: tone = `NM8 << 1;
        13'd2039: tone = `NM8 << 1;
        13'd2040: tone = `NM2 << 2;
        13'd2041: tone = `NM2 << 2;
        13'd2042: tone = `NM2 << 2;
        13'd2043: tone = `NM2 << 2;
        13'd2044: tone = `NM2 <<2;
        13'd2045: tone = `NM2 << 2;
        13'd2046: tone = `NM2 << 2;
        13'd2047: tone = `NM2 << 2;
        
        13'd2048: tone = `NM2 << 2;
        13'd2049: tone = `NM2 << 2;
        13'd2050: tone = `NM2 << 2;
        13'd2051: tone = `NM2 << 2;
        13'd2052: tone = `NM2 << 2;
        13'd2053: tone = `NM2 << 2;
        13'd2054: tone = `NM2 << 2;
        13'd2055: tone = `NM2 << 2;
        13'd2056: tone = `NM1 << 2;
        13'd2057: tone = `NM1 << 2;
        13'd2058: tone = `NM1 << 2;
        13'd2059: tone = `NM1 << 2;
        13'd2060: tone = `NM1 << 2;
        13'd2061: tone = `NM1 << 2;
        13'd2062: tone = `NM1 << 2;
        13'd2063: tone = `NM1 << 2;
        
        13'd2064: tone = `NM11 <<1;
        13'd2065: tone = `NM11 <<1;
        13'd2066: tone = `NM11 <<1;
        13'd2067: tone = `NM11 <<1;
        13'd2068: tone = `NM11 <<1;
        13'd2069: tone = `NM11 <<1;
        13'd2070: tone = `NM11 <<1;
        13'd2071: tone = `NM0;
        13'd2072: tone = `NM11 <<1;
        13'd2073: tone = `NM11 <<1;
        13'd2074: tone = `NM11 <<1;
        13'd2075: tone = `NM11 <<1;
        13'd2076: tone = `NM11 <<1;
        13'd2077: tone = `NM11 <<1;
        13'd2078: tone = `NM11 <<1;
        13'd2079: tone = `NM11 <<1;
        
        13'd2080: tone = `NM11 <<1;
        13'd2081: tone = `NM11 <<1;
        13'd2082: tone = `NM11 <<1;
        13'd2083: tone = `NM11 <<1;
        13'd2084: tone = `NM11 <<1;
        13'd2085: tone = `NM11 <<1;
        13'd2086: tone = `NM11 <<1;
        13'd2087: tone = `NM0;
        13'd2088: tone = `NM11 <<1;
        13'd2089: tone = `NM11 <<1;
        13'd2090: tone = `NM11 <<1;
        13'd2091: tone = `NM11 <<1;
        13'd2092: tone = `NM11 <<1;
        13'd2093: tone = `NM11 <<1;
        13'd2094: tone = `NM11 <<1;
        13'd2095: tone = `NM11 <<1;
        
        13'd2096: tone = `NM1 <<2;
        13'd2097: tone = `NM1 <<2;
        13'd2098: tone = `NM1 <<2;
        13'd2099: tone = `NM1 <<2;
        13'd2100: tone = `NM1 <<2;
        13'd2101: tone = `NM1 <<2;
        13'd2102: tone = `NM1 <<2;
        13'd2103: tone = `NM1 <<2;
        13'd2104: tone = `NM6 << 1;
        13'd2105: tone = `NM6 << 1;
        13'd2106: tone = `NM6 << 1;
        13'd2107: tone = `NM6 << 1;
        13'd2108: tone = `NM6 << 1;
        13'd2109: tone = `NM6 << 1;
        13'd2110: tone = `NM6 << 1;
        13'd2111: tone = `NM6 << 1;
        
        13'd2112: tone = `NM8 << 1;
        13'd2113: tone = `NM8 << 1;
        13'd2114: tone = `NM8 << 1;
        13'd2115: tone = `NM8 << 1;
        13'd2116: tone = `NM8 << 1;
        13'd2117: tone = `NM8 << 1;
        13'd2118: tone = `NM8 << 1;
        13'd2119: tone = `NM8 << 1;
        13'd2120: tone = `NM8 << 1;
        13'd2121: tone = `NM8 << 1;
        13'd2122: tone = `NM8 << 1;
        13'd2123: tone = `NM8 << 1;
        13'd2124: tone = `NM8 << 1;
        13'd2125: tone = `NM8 << 1;
        13'd2126: tone = `NM8 << 1;
        13'd2127: tone = `NM8 << 1;
        
        13'd2128: tone = `NM0;
        13'd2129: tone = `NM0;
        13'd2130: tone = `NM0;
        13'd2131: tone = `NM0;
        13'd2132: tone = `NM0;
        13'd2133: tone = `NM0;
        13'd2134: tone = `NM0;
        13'd2135: tone = `NM0;
        13'd2136: tone = `NM8 << 1;
        13'd2137: tone = `NM8 << 1;
        13'd2138: tone = `NM8 << 1;
        13'd2139: tone = `NM8 << 1;
        13'd2140: tone = `NM8 << 1;
        13'd2141: tone = `NM8 << 1;
        13'd2142: tone = `NM8 << 1;
        13'd2143: tone = `NM8 << 1;
        
        13'd2144: tone = `NM11 << 1;
        13'd2145: tone = `NM11 << 1;
        13'd2146: tone = `NM11 << 1;
        13'd2147: tone = `NM11 << 1;
        13'd2148: tone = `NM11 << 1;
        13'd2149: tone = `NM11 << 1;
        13'd2150: tone = `NM11 << 1;
        13'd2151: tone = `NM0;
        13'd2152: tone = `NM11 << 1;
        13'd2153: tone = `NM11 << 1;
        13'd2154: tone = `NM11 << 1;
        13'd2155: tone = `NM11 << 1;
        13'd2156: tone = `NM11 << 1;
        13'd2157: tone = `NM11 << 1;
        13'd2158: tone = `NM11 << 1;
        13'd2159: tone = `NM11 << 1;
        
        13'd2160: tone = `NM0;
        13'd2161: tone = `NM0;
        13'd2162: tone = `NM0;
        13'd2163: tone = `NM0;
        13'd2164: tone = `NM0;
        13'd2165: tone = `NM0;
        13'd2166: tone = `NM0;
        13'd2167: tone = `NM0;
        13'd2168: tone = `NM2 << 2;
        13'd2169: tone = `NM2 << 2;
        13'd2170: tone = `NM2 << 2;
        13'd2171: tone = `NM2 << 2;
        13'd2172: tone = `NM2 << 2;
        13'd2173: tone = `NM2 << 2;
        13'd2174: tone = `NM2 << 2;
        13'd2175: tone = `NM2 << 2;
        
        13'd2176: tone = `NM2 << 2;
        13'd2177: tone = `NM2 << 2;
        13'd2178: tone = `NM2 << 2;
        13'd2179: tone = `NM2 << 2;
        13'd2180: tone = `NM2 << 2;
        13'd2181: tone = `NM2 << 2;
        13'd2182: tone = `NM2 << 2;
        13'd2183: tone = `NM2 << 2;
        13'd2184: tone = `NM1 << 2;
        13'd2185: tone = `NM1 << 2;
        13'd2186: tone = `NM1 << 2;
        13'd2187: tone = `NM1 << 2;
        13'd2188: tone = `NM1 << 2;
        13'd2189: tone = `NM1 << 2;
        13'd2190: tone = `NM1 << 2;
        13'd2191: tone = `NM1 << 2;
        
        13'd2192: tone = `NM11 << 1;
        13'd2193: tone = `NM11 << 1;
        13'd2194: tone = `NM11 << 1;
        13'd2195: tone = `NM11 << 1;
        13'd2196: tone = `NM11 << 1;
        13'd2197: tone = `NM11 << 1;
        13'd2198: tone = `NM11 << 1;
        13'd2199: tone = `NM0;
        13'd2200: tone = `NM11 << 1;
        13'd2201: tone = `NM11 << 1;
        13'd2202: tone = `NM11 << 1;
        13'd2203: tone = `NM11 << 1;
        13'd2204: tone = `NM11 << 1;
        13'd2205: tone = `NM11 << 1;
        13'd2206: tone = `NM11 << 1;
        13'd2207: tone = `NM11 << 1;
        
        13'd2208: tone = `NM11 << 1;
        13'd2209: tone = `NM11 << 1;
        13'd2210: tone = `NM11 << 1;
        13'd2211: tone = `NM11 << 1;
        13'd2212: tone = `NM11 << 1;
        13'd2213: tone = `NM11 << 1;
        13'd2214: tone = `NM11 << 1;
        13'd2215: tone = `NM0;
        13'd2216: tone = `NM11 << 1;
        13'd2217: tone = `NM11 << 1;
        13'd2218: tone = `NM11 << 1;
        13'd2219: tone = `NM11 << 1;
        13'd2220: tone = `NM11 << 1;
        13'd2221: tone = `NM11 << 1;
        13'd2222: tone = `NM11 << 1;
        13'd2223: tone = `NM11 << 1;
        
        13'd2224: tone = `NM1 <<2;
        13'd2225: tone = `NM1 <<2;
        13'd2226: tone = `NM1 <<2;
        13'd2227: tone = `NM1 <<2;
        13'd2228: tone = `NM1 <<2;
        13'd2229: tone = `NM1 <<2;
        13'd2230: tone = `NM1 <<2;
        13'd2231: tone = `NM1 <<2;
        13'd2232: tone = `NM6 << 1;
        13'd2233: tone = `NM6 << 1;
        13'd2234: tone = `NM6 << 1;
        13'd2235: tone = `NM6 << 1;
        13'd2236: tone = `NM6 << 1;
        13'd2237: tone = `NM6 << 1;
        13'd2238: tone = `NM6 << 1;
        13'd2239: tone = `NM6 << 1;
        
        13'd2240: tone = `NM8 << 1;
        13'd2241: tone = `NM8 << 1;
        13'd2242: tone = `NM8 << 1;
        13'd2243: tone = `NM8 << 1;
        13'd2244: tone = `NM8 << 1;
        13'd2245: tone = `NM8 << 1;
        13'd2246: tone = `NM8 << 1;
        13'd2247: tone = `NM8 << 1;
        13'd2248: tone = `NM8 << 1;
        13'd2249: tone = `NM8 << 1;
        13'd2250: tone = `NM8 << 1;
        13'd2251: tone = `NM8 << 1;
        13'd2252: tone = `NM8 << 1;
        13'd2253: tone = `NM8 << 1;
        13'd2254: tone = `NM8 << 1;
        13'd2255: tone = `NM8 << 1;
        
        13'd2256: tone = `NM0;
        13'd2257: tone = `NM0;
        13'd2258: tone = `NM0;
        13'd2259: tone = `NM0;
        13'd2260: tone = `NM0;
        13'd2261: tone = `NM0;
        13'd2262: tone = `NM0;
        13'd2263: tone = `NM0;
        13'd2264: tone = `NM8 << 1;
        13'd2265: tone = `NM8 << 1;
        13'd2266: tone = `NM8 << 1;
        13'd2267: tone = `NM8 << 1;
        13'd2268: tone = `NM8 << 1;
        13'd2269: tone = `NM8 << 1;
        13'd2270: tone = `NM8 << 1;
        13'd2271: tone = `NM8 << 1;
        
        13'd2272: tone = `NM11 << 1;
        13'd2273: tone = `NM11 << 1;
        13'd2274: tone = `NM11 << 1;
        13'd2275: tone = `NM11 << 1;
        13'd2276: tone = `NM11 << 1;
        13'd2277: tone = `NM11 << 1;
        13'd2278: tone = `NM11 << 1;
        13'd2279: tone = `NM0;
        13'd2280: tone = `NM11 << 1;
        13'd2281: tone = `NM11 << 1;
        13'd2282: tone = `NM11 << 1;
        13'd2283: tone = `NM11 << 1;
        13'd2284: tone = `NM11 << 1;
        13'd2285: tone = `NM11 << 1;
        13'd2286: tone = `NM11 << 1;
        13'd2287: tone = `NM11 << 1;
        
        13'd2288: tone = `NM8 << 1;
        13'd2289: tone = `NM8 << 1;
        13'd2290: tone = `NM8 << 1;
        13'd2291: tone = `NM8 << 1;
        13'd2292: tone = `NM8 << 1;
        13'd2293: tone = `NM8 << 1;
        13'd2294: tone = `NM8 << 1;
        13'd2295: tone = `NM8 << 1;
        13'd2296: tone = `NM2 << 2;
        13'd2297: tone = `NM2 << 2;
        13'd2298: tone = `NM2 << 2;
        13'd2299: tone = `NM2 << 2;
        13'd2300: tone = `NM2 << 2;
        13'd2301: tone = `NM2 << 2;
        13'd2302: tone = `NM2 << 2;
        13'd2303: tone = `NM2 << 2;
        
        13'd2304: tone = `NM2 << 2;
        13'd2305: tone = `NM2 << 2;
        13'd2306: tone = `NM2 << 2;
        13'd2307: tone = `NM2 << 2;
        13'd2308: tone = `NM2 << 2;
        13'd2309: tone = `NM2 << 2;
        13'd2310: tone = `NM2 << 2;
        13'd2311: tone = `NM2 << 2;
        13'd2312: tone = `NM1 << 2;
        13'd2313: tone = `NM1 << 2;
        13'd2314: tone = `NM1 << 2;
        13'd2315: tone = `NM1 << 2;
        13'd2316: tone = `NM1 << 2;
        13'd2317: tone = `NM1 << 2;
        13'd2318: tone = `NM1 << 2;
        13'd2319: tone = `NM1 << 2;
        
        13'd2320: tone = `NM11 << 1;
        13'd2321: tone = `NM11 << 1;
        13'd2322: tone = `NM11 << 1;
        13'd2323: tone = `NM11 << 1;
        13'd2324: tone = `NM11 << 1;
        13'd2325: tone = `NM11 << 1;
        13'd2326: tone = `NM11 << 1;
        13'd2327: tone = `NM0;
        13'd2328: tone = `NM11 << 1;
        13'd2329: tone = `NM11 << 1;
        13'd2330: tone = `NM11 << 1;
        13'd2331: tone = `NM11 << 1;
        13'd2332: tone = `NM11 << 1;
        13'd2333: tone = `NM11 << 1;
        13'd2334: tone = `NM11 << 1;
        13'd2335: tone = `NM11 << 1;
        
        13'd2336: tone = `NM11 << 1;
        13'd2337: tone = `NM11 << 1;
        13'd2338: tone = `NM11 << 1;
        13'd2339: tone = `NM11 << 1;
        13'd2340: tone = `NM11 << 1;
        13'd2341: tone = `NM11 << 1;
        13'd2342: tone = `NM11 << 1;
        13'd2343: tone = `NM0;
        13'd2344: tone = `NM11 << 1;
        13'd2345: tone = `NM11 << 1;
        13'd2346: tone = `NM11 << 1;
        13'd2347: tone = `NM11 << 1;
        13'd2348: tone = `NM11 << 1;
        13'd2349: tone = `NM11 << 1;
        13'd2350: tone = `NM11 << 1;
        13'd2351: tone = `NM11 << 1;
        
        13'd2352: tone = `NM1 << 2;
        13'd2353: tone = `NM1 << 2;
        13'd2354: tone = `NM1 << 2;
        13'd2355: tone = `NM1 << 2;
        13'd2356: tone = `NM1 << 2;
        13'd2357: tone = `NM1 << 2;
        13'd2358: tone = `NM1 << 2;
        13'd2359: tone = `NM1 << 2;
        13'd2360: tone = `NM6 << 1;
        13'd2361: tone = `NM6 << 1;
        13'd2362: tone = `NM6 << 1;
        13'd2363: tone = `NM6 << 1;
        13'd2364: tone = `NM6 << 1;
        13'd2365: tone = `NM6 << 1;
        13'd2366: tone = `NM6 << 1;
        13'd2367: tone = `NM6 << 1;
        
        13'd2368: tone = `NM8 << 1;
        13'd2369: tone = `NM8 << 1;
        13'd2370: tone = `NM8 << 1;
        13'd2371: tone = `NM8 << 1;
        13'd2372: tone = `NM8 << 1;
        13'd2373: tone = `NM8 << 1;
        13'd2374: tone = `NM8 << 1;
        13'd2375: tone = `NM8 << 1;
        13'd2376: tone = `NM8 << 1;
        13'd2377: tone = `NM8 << 1;
        13'd2378: tone = `NM8 << 1;
        13'd2379: tone = `NM8 << 1;
        13'd2380: tone = `NM8 << 1;
        13'd2381: tone = `NM8 << 1;
        13'd2382: tone = `NM8 << 1;
        13'd2383: tone = `NM0;
        
        13'd2384: tone = `NM8 << 1;
        13'd2385: tone = `NM8 << 1;
        13'd2386: tone = `NM8 << 1;
        13'd2387: tone = `NM8 << 1;
        13'd2388: tone = `NM8 << 1;
        13'd2389: tone = `NM8 << 1;
        13'd2390: tone = `NM8 << 1;
        13'd2391: tone = `NM8 << 1;
        13'd2392: tone = `NM10 << 1;
        13'd2393: tone = `NM10 << 1;
        13'd2394: tone = `NM10 << 1;
        13'd2395: tone = `NM10 << 1;
        13'd2396: tone = `NM10 << 1;
        13'd2397: tone = `NM10 << 1;
        13'd2398: tone = `NM10 << 1;
        13'd2399: tone = `NM10 << 1;
        
        13'd2400: tone = `NM11 << 1;
        13'd2401: tone = `NM11 << 1;
        13'd2402: tone = `NM11 << 1;
        13'd2403: tone = `NM11 << 1;
        13'd2404: tone = `NM11 << 1;
        13'd2405: tone = `NM11 << 1;
        13'd2406: tone = `NM11 << 1;
        13'd2407: tone = `NM11 << 1;
        13'd2408: tone = `NM10 << 1;
        13'd2409: tone = `NM10 << 1;
        13'd2410: tone = `NM10 << 1;
        13'd2411: tone = `NM10 << 1;
        13'd2412: tone = `NM10 << 1;
        13'd2413: tone = `NM10 << 1;
        13'd2414: tone = `NM10 << 1;
        13'd2415: tone = `NM10 << 1;
        
        13'd2416: tone = `NM8 << 1;
        13'd2417: tone = `NM8 << 1;
        13'd2418: tone = `NM8 << 1;
        13'd2419: tone = `NM8 << 1;
        13'd2420: tone = `NM8 << 1;
        13'd2421: tone = `NM8 << 1;
        13'd2422: tone = `NM8 << 1;
        13'd2423: tone = `NM0;
        13'd2424: tone = `NM8 << 1;
        13'd2425: tone = `NM8 << 1;
        13'd2426: tone = `NM8 << 1;
        13'd2427: tone = `NM8 << 1;
        13'd2428: tone = `NM8 << 1;
        13'd2429: tone = `NM8 << 1;
        13'd2430: tone = `NM8 << 1;
        13'd2431: tone = `NM8 << 1;
        
        13'd2432: tone = `NM8 << 1;
        13'd2433: tone = `NM8 << 1;
        13'd2434: tone = `NM8 << 1;
        13'd2435: tone = `NM8 << 1;
        13'd2436: tone = `NM8 << 1;
        13'd2437: tone = `NM8 << 1;
        13'd2438: tone = `NM8 << 1;
        13'd2439: tone = `NM8 << 1;
        13'd2440: tone = `NM8 << 1;
        13'd2441: tone = `NM8 << 1;
        13'd2442: tone = `NM8 << 1;
        13'd2443: tone = `NM8 << 1;
        13'd2444: tone = `NM8 << 1;
        13'd2445: tone = `NM8 << 1;
        13'd2446: tone = `NM8 << 1;
        13'd2447: tone = `NM8 << 1;
        
        13'd2448: tone = `NM0;
        13'd2449: tone = `NM0;
        13'd2450: tone = `NM0;
        13'd2451: tone = `NM0;
        13'd2452: tone = `NM0;
        13'd2453: tone = `NM0;
        13'd2454: tone = `NM0;
        13'd2455: tone = `NM0;
        13'd2456: tone = `NM8 << 1;
        13'd2457: tone = `NM8 << 1;
        13'd2458: tone = `NM8 << 1;
        13'd2459: tone = `NM8 << 1;
        13'd2460: tone = `NM8 << 1;
        13'd2461: tone = `NM8 << 1;
        13'd2462: tone = `NM8 << 1;
        13'd2463: tone = `NM8 << 1;
        
        13'd2464: tone = `NM8 << 1;
        13'd2465: tone = `NM8 << 1;
        13'd2466: tone = `NM8 << 1;
        13'd2467: tone = `NM8 << 1;
        13'd2468: tone = `NM8 << 1;
        13'd2469: tone = `NM8 << 1;
        13'd2470: tone = `NM8 << 1;
        13'd2471: tone = `NM8 << 1;
        13'd2472: tone = `NM8 << 1;
        13'd2473: tone = `NM8 << 1;
        13'd2474: tone = `NM8 << 1;
        13'd2475: tone = `NM8 << 1;
        13'd2476: tone = `NM8 << 1;
        13'd2477: tone = `NM8 << 1;
        13'd2478: tone = `NM8 << 1;
        13'd2479: tone = `NM8 << 1;
        
        13'd2480: tone = `NM0;
        13'd2481: tone = `NM0;
        13'd2482: tone = `NM0;
        13'd2483: tone = `NM0;
        13'd2484: tone = `NM0;
        13'd2485: tone = `NM0;
        13'd2486: tone = `NM0;
        13'd2487: tone = `NM0;
        13'd2488: tone = `NM8 << 1;
        13'd2489: tone = `NM8 << 1;
        13'd2490: tone = `NM8 << 1;
        13'd2491: tone = `NM8 << 1;
        13'd2492: tone = `NM8 << 1;
        13'd2493: tone = `NM8 << 1;
        13'd2494: tone = `NM8 << 1;
        13'd2495: tone = `NM8 << 1;
        13'd2496: tone = `NM8 << 1;

        13'd2497: tone = `NM8 << 1;
        13'd2498: tone = `NM8 << 1;
        13'd2499: tone = `NM8 << 1;
        13'd2500: tone = `NM8 << 1;
        13'd2501: tone = `NM8 << 1;
        13'd2502: tone = `NM8 << 1;
        13'd2503: tone = `NM8 << 1;
        13'd2504: tone = `NM8 << 1;
        13'd2505: tone = `NM8 << 1;
        13'd2506: tone = `NM8 << 1;
        13'd2507: tone = `NM8 << 1;
        13'd2508: tone = `NM8 << 1;
        13'd2509: tone = `NM8 << 1;
        13'd2510: tone = `NM8 << 1;
        13'd2511: tone = `NM8 << 1;
        13'd2512: tone = `NM8 << 1;
        
        13'd2513: tone = `NM8 << 1;
        13'd2514: tone = `NM8 << 1;
        13'd2515: tone = `NM8 << 1;
        13'd2516: tone = `NM8 << 1;
        13'd2517: tone = `NM8 << 1;
        13'd2518: tone = `NM8 << 1;
        13'd2519: tone = `NM8 << 1;
        13'd2520: tone = `NM8 << 1;
        13'd2521: tone = `NM8 << 1;
        13'd2522: tone = `NM8 << 1;
        13'd2523: tone = `NM8 << 1;
        13'd2524: tone = `NM8 << 1;
        13'd2525: tone = `NM8 << 1;
        13'd2526: tone = `NM8 << 1;
        13'd2527: tone = `NM8 << 1;
        
        13'd2528: tone = `NM0;
        13'd2529: tone = `NM0;
        13'd2530: tone = `NM0;
        13'd2531: tone = `NM0;
        13'd2532: tone = `NM0;
        13'd2533: tone = `NM0;
        13'd2534: tone = `NM0;
        13'd2535: tone = `NM0;
        13'd2536: tone = `NM11 << 1;
        13'd2537: tone = `NM11 << 1;
        13'd2538: tone = `NM11 << 1;
        13'd2539: tone = `NM11 << 1;
        13'd2540: tone = `NM11 << 1;
        13'd2541: tone = `NM11 << 1;
        13'd2542: tone = `NM11 << 1;
        13'd2543: tone = `NM0;
        
        13'd2544: tone = `NM11 << 1;
        13'd2545: tone = `NM11 << 1;
        13'd2546: tone = `NM11 << 1;
        13'd2547: tone = `NM11 << 1;
        13'd2548: tone = `NM11 << 1;
        13'd2549: tone = `NM11 << 1;
        13'd2550: tone = `NM11 << 1;
        13'd2551: tone = `NM0;
        13'd2552: tone = `NM8 << 1;
        13'd2553: tone = `NM8 << 1;
        13'd2554: tone = `NM8 << 1;
        13'd2555: tone = `NM8 << 1;
        13'd2556: tone = `NM8 << 1;
        13'd2557: tone = `NM8 << 1;
        13'd2558: tone = `NM8 << 1;
        13'd2559: tone = `NM0;
        
        13'd2560: tone = `NM11 << 1;
        13'd2561: tone = `NM11 << 1;
        13'd2562: tone = `NM11 << 1;
        13'd2563: tone = `NM11 << 1;
        13'd2564: tone = `NM11 << 1;
        13'd2565: tone = `NM11 << 1;
        13'd2566: tone = `NM11 << 1;
        13'd2567: tone = `NM11 << 1;
        13'd2568: tone = `NM8 << 1;
        13'd2569: tone = `NM8 << 1;
        13'd2570: tone = `NM8 << 1;
        13'd2571: tone = `NM8 << 1;
        13'd2572: tone = `NM8 << 1;
        13'd2573: tone = `NM8 << 1;
        13'd2574: tone = `NM8 << 1;
        13'd2575: tone = `NM8 << 1;
        
        13'd2576: tone = `NM11 << 1;
        13'd2577: tone = `NM11 << 1;
        13'd2578: tone = `NM11 << 1;
        13'd2579: tone = `NM11 << 1;
        13'd2580: tone = `NM11 << 1;
        13'd2581: tone = `NM11 << 1;
        13'd2582: tone = `NM11 << 1;
        13'd2583: tone = `NM11 << 1;
        13'd2584: tone = `NM11 << 1;
        13'd2585: tone = `NM11 << 1;
        13'd2586: tone = `NM11 << 1;
        13'd2587: tone = `NM11 << 1;
        13'd2588: tone = `NM0;
        13'd2589: tone = `NM0;
        13'd2590: tone = `NM0;
        13'd2591: tone = `NM0;
        
        13'd2592: tone = `NM11 << 1;
        13'd2593: tone = `NM11 << 1;
        13'd2594: tone = `NM11 << 1;
        13'd2595: tone = `NM11 << 1;
        13'd2596: tone = `NM11 << 1;
        13'd2597: tone = `NM11 << 1;
        13'd2598: tone = `NM11 << 1;
        13'd2599: tone = `NM11 << 1;
        13'd2600: tone = `NM11 << 1;
        13'd2601: tone = `NM11 << 1;
        13'd2602: tone = `NM11 << 1;
        13'd2603: tone = `NM11 << 1;
        13'd2604: tone = `NM11 << 1;
        13'd2605: tone = `NM11 << 1;
        13'd2606: tone = `NM11 << 1;
        13'd2607: tone = `NM0;
        
        13'd2608: tone = `NM11 << 1;
        13'd2609: tone = `NM11 << 1;
        13'd2610: tone = `NM11 << 1;
        13'd2611: tone = `NM11 << 1;
        13'd2612: tone = `NM11 << 1;
        13'd2613: tone = `NM11 << 1;
        13'd2614: tone = `NM11 << 1;
        13'd2615: tone = `NM0;
        13'd2616: tone = `NM11 << 1;
        13'd2617: tone = `NM11 << 1;
        13'd2618: tone = `NM11 << 1;
        13'd2619: tone = `NM11 << 1;
        13'd2620: tone = `NM11 << 1;
        13'd2621: tone = `NM11 << 1;
        13'd2622: tone = `NM11 << 1;
        13'd2623: tone = `NM0;
        
        13'd2624: tone = `NM11 << 1;
        13'd2625: tone = `NM11 << 1;
        13'd2626: tone = `NM11 << 1;
        13'd2627: tone = `NM11 << 1;
        13'd2628: tone = `NM11 << 1;
        13'd2629: tone = `NM11 << 1;
        13'd2630: tone = `NM11 << 1;
        13'd2631: tone = `NM11 << 1;
        13'd2632: tone = `NM10 << 1;
        13'd2633: tone = `NM10 << 1;
        13'd2634: tone = `NM10 << 1;
        13'd2635: tone = `NM10 << 1;
        13'd2636: tone = `NM10 << 1;
        13'd2637: tone = `NM10 << 1;
        13'd2638: tone = `NM10 << 1;
        13'd2639: tone = `NM10 << 1;
        
        13'd2640: tone = `NM8 << 1;
        13'd2641: tone = `NM8 << 1;
        13'd2642: tone = `NM8 << 1;
        13'd2643: tone = `NM8 << 1;
        13'd2644: tone = `NM8 << 1;
        13'd2645: tone = `NM8 << 1;
        13'd2646: tone = `NM8 << 1;
        13'd2647: tone = `NM0;
        13'd2648: tone = `NM8 << 1;
        13'd2649: tone = `NM8 << 1;
        13'd2650: tone = `NM8 << 1;
        13'd2651: tone = `NM8 << 1;
        13'd2652: tone = `NM8 <<1;
        13'd2653: tone = `NM8 << 1;
        13'd2654: tone = `NM8 << 1;
        13'd2655: tone = `NM0;
        
        13'd2656: tone = `NM0;
        13'd2657: tone = `NM0;
        13'd2658: tone = `NM0;
        13'd2659: tone = `NM0;
        13'd2660: tone = `NM0;
        13'd2661: tone = `NM0;
        13'd2662: tone = `NM0;
        13'd2663: tone = `NM0;
        13'd2664: tone = `NM11 << 1;
        13'd2665: tone = `NM11 << 1;
        13'd2666: tone = `NM11 << 1;
        13'd2667: tone = `NM11 << 1;
        13'd2668: tone = `NM11 << 1;
        13'd2669: tone = `NM11 << 1;
        13'd2670: tone = `NM11 << 1;
        13'd2671: tone = `NM0;
        
        13'd2672: tone = `NM11 << 1;
        13'd2673: tone = `NM11 << 1;
        13'd2674: tone = `NM11 << 1;
        13'd2675: tone = `NM11 << 1;
        13'd2676: tone = `NM11 << 1;
        13'd2677: tone = `NM11 << 1;
        13'd2678: tone = `NM11 << 1;
        13'd2679: tone = `NM11 << 1;
        13'd2680: tone = `NM8 << 1;
        13'd2681: tone = `NM8 << 1;
        13'd2682: tone = `NM8 << 1;
        13'd2683: tone = `NM8 << 1;
        13'd2684: tone = `NM8 << 1;
        13'd2685: tone = `NM8 << 1;
        13'd2686: tone = `NM8 << 1;
        13'd2687: tone = `NM8 << 1;
        
        13'd2688: tone = `NM11 << 1;
        13'd2689: tone = `NM11 << 1;
        13'd2690: tone = `NM11 << 1;
        13'd2691: tone = `NM11 << 1;
        13'd2692: tone = `NM11 << 1;
        13'd2693: tone = `NM11 << 1;
        13'd2694: tone = `NM11 << 1;
        13'd2695: tone = `NM11 << 1;
        13'd2696: tone = `NM8 << 1;
        13'd2697: tone = `NM8 << 1;
        13'd2698: tone = `NM8 << 1;
        13'd2699: tone = `NM8 << 1;
        13'd2700: tone = `NM8 << 1;
        13'd2701: tone = `NM8 << 1;
        13'd2702: tone = `NM8 << 1;
        13'd2703: tone = `NM8 << 1;
        
        13'd2704: tone = `NM11 << 1;
        13'd2705: tone = `NM11 << 1;
        13'd2706: tone = `NM11 << 1;
        13'd2707: tone = `NM11 << 1;
        13'd2708: tone = `NM11 << 1;
        13'd2709: tone = `NM11 << 1;
        13'd2710: tone = `NM11 << 1;
        13'd2711: tone = `NM11 << 1;
        13'd2712: tone = `NM11 << 1;
        13'd2713: tone = `NM11 << 1;
        13'd2714: tone = `NM11 << 1;
        13'd2715: tone = `NM11 << 1;
        13'd2716: tone = `NM0;
        13'd2717: tone = `NM0;
        13'd2718: tone = `NM0;
        13'd2719: tone = `NM0;
        
        13'd2720: tone = `NM11 << 1;
        13'd2721: tone = `NM11 << 1;
        13'd2722: tone = `NM11 << 1;
        13'd2723: tone = `NM11 << 1;
        13'd2724: tone = `NM11 << 1;
        13'd2725: tone = `NM11 << 1;
        13'd2726: tone = `NM11 << 1;
        13'd2727: tone = `NM11 << 1;
        13'd2728: tone = `NM11 << 1;
        13'd2729: tone = `NM11 << 1;
        13'd2730: tone = `NM11 << 1;
        13'd2731: tone = `NM11 << 1;
        13'd2732: tone = `NM11 << 1;
        13'd2733: tone = `NM11 << 1;
        13'd2734: tone = `NM11 << 1;
        13'd2735: tone = `NM0;
        
        13'd2736: tone = `NM11 << 1;
        13'd2737: tone = `NM11 << 1;
        13'd2738: tone = `NM11 << 1;
        13'd2739: tone = `NM11 << 1;
        13'd2740: tone = `NM11 << 1;
        13'd2741: tone = `NM11 << 1;
        13'd2742: tone = `NM11 << 1;
        13'd2743: tone = `NM0;
        13'd2744: tone = `NM11 << 1;
        13'd2745: tone = `NM11 << 1;
        13'd2746: tone = `NM11 << 1;
        13'd2747: tone = `NM11 << 1;
        13'd2748: tone = `NM11 << 1;
        13'd2749: tone = `NM11 << 1;
        13'd2750: tone = `NM11 << 1;
        13'd2751: tone = `NM0;
        
        13'd2752: tone = `NM1 << 2;
        13'd2753: tone = `NM1 << 2;
        13'd2754: tone = `NM1 << 2;
        13'd2755: tone = `NM1 << 2;
        13'd2756: tone = `NM1 << 2;
        13'd2757: tone = `NM1 << 2;
        13'd2758: tone = `NM1 << 2;
        13'd2759: tone = `NM1 << 2;
        13'd2760: tone = `NM11 << 1;
        13'd2761: tone = `NM11 << 1;
        13'd2762: tone = `NM11 << 1;
        13'd2763: tone = `NM11 << 1;
        13'd2764: tone = `NM11 << 1;
        13'd2765: tone = `NM11 << 1;
        13'd2766: tone = `NM11 << 1;
        13'd2767: tone = `NM11 << 1;
        
        13'd2768: tone = `NM8 << 1;
        13'd2769: tone = `NM8 << 1;
        13'd2770: tone = `NM8 << 1;
        13'd2771: tone = `NM8 << 1;
        13'd2772: tone = `NM8 << 1;
        13'd2773: tone = `NM8 << 1;
        13'd2774: tone = `NM8 << 1;
        13'd2775: tone = `NM0;
        13'd2776: tone = `NM8 << 1;
        13'd2777: tone = `NM8 << 1;
        13'd2778: tone = `NM8 << 1;
        13'd2779: tone = `NM8 << 1;
        13'd2780: tone = `NM8 << 1;
        13'd2781: tone = `NM8 << 1;
        13'd2782: tone = `NM8 << 1;
        13'd2783: tone = `NM8 << 1;
        
        13'd2784: tone = `NM0;
        13'd2785: tone = `NM0;
        13'd2786: tone = `NM0;
        13'd2787: tone = `NM0;
        13'd2788: tone = `NM0;
        13'd2789: tone = `NM0;
        13'd2790: tone = `NM0;
        13'd2791: tone = `NM0;
        13'd2792: tone = `NM11 << 1;
        13'd2793: tone = `NM11 << 1;
        13'd2794: tone = `NM11 << 1;
        13'd2795: tone = `NM11 << 1;
        13'd2796: tone = `NM11 << 1;
        13'd2797: tone = `NM11 << 1;
        13'd2798: tone = `NM11 << 1;
        13'd2799: tone = `NM0;
        
        13'd2800: tone = `NM11 << 1;
        13'd2801: tone = `NM11 << 1;
        13'd2802: tone = `NM11 << 1;
        13'd2803: tone = `NM11 << 1;
        13'd2804: tone = `NM11 << 1;
        13'd2805: tone = `NM11 << 1;
        13'd2806: tone = `NM11 << 1;
        13'd2807: tone = `NM0;
        13'd2808: tone = `NM8 << 1;
        13'd2809: tone = `NM8 << 1;
        13'd2810: tone = `NM8 << 1;
        13'd2811: tone = `NM8 << 1;
        13'd2812: tone = `NM8 << 1;
        13'd2813: tone = `NM8 << 1;
        13'd2814: tone = `NM8 << 1;
        13'd2815: tone = `NM8 << 1;
        
        13'd2816: tone = `NM11 << 1;
        13'd2817: tone = `NM11 << 1;
        13'd2818: tone = `NM11 << 1;
        13'd2819: tone = `NM11 << 1;
        13'd2820: tone = `NM11 << 1;
        13'd2821: tone = `NM11 << 1;
        13'd2822: tone = `NM11 << 1;
        13'd2823: tone = `NM11 << 1;
        13'd2824: tone = `NM8 << 1;
        13'd2825: tone = `NM8 << 1;
        13'd2826: tone = `NM8 << 1;
        13'd2827: tone = `NM8 << 1;
        13'd2828: tone = `NM8 << 1;
        13'd2829: tone = `NM8 << 1;
        13'd2830: tone = `NM8 << 1;
        13'd2831: tone = `NM8 << 1;
        
        13'd2832: tone = `NM11 << 1;
        13'd2833: tone = `NM11 << 1;
        13'd2834: tone = `NM11 << 1;
        13'd2835: tone = `NM11 << 1;
        13'd2836: tone = `NM11 << 1;
        13'd2837: tone = `NM11 << 1;
        13'd2838: tone = `NM11 << 1;
        13'd2839: tone = `NM11 << 1;
        13'd2840: tone = `NM11 << 1;
        13'd2841: tone = `NM11 << 1;
        13'd2842: tone = `NM11 << 1;
        13'd2843: tone = `NM11 << 1;
        13'd2844: tone = `NM0;
        13'd2845: tone = `NM0;
        13'd2846: tone = `NM0;
        13'd2847: tone = `NM0;
        
        13'd2848: tone = `NM11 << 1;
        13'd2849: tone = `NM11 << 1;
        13'd2850: tone = `NM11 << 1;
        13'd2851: tone = `NM11 << 1;
        13'd2852: tone = `NM11 << 1;
        13'd2853: tone = `NM11 << 1;
        13'd2854: tone = `NM11 << 1;
        13'd2855: tone = `NM11 << 1;
        13'd2856: tone = `NM11 << 1;
        13'd2857: tone = `NM11 << 1;
        13'd2858: tone = `NM11 << 1;
        13'd2859: tone = `NM11 << 1;
        13'd2860: tone = `NM11 << 1;
        13'd2861: tone = `NM11 << 1;
        13'd2862: tone = `NM11 << 1;
        13'd2863: tone = `NM0;
        
        13'd2864: tone = `NM11 << 1;
        13'd2865: tone = `NM11 << 1;
        13'd2866: tone = `NM11 << 1;
        13'd2867: tone = `NM11 << 1;
        13'd2868: tone = `NM11 << 1;
        13'd2869: tone = `NM11 << 1;
        13'd2870: tone = `NM11 << 1;
        13'd2871: tone = `NM0;
        13'd2872: tone = `NM11 << 1;
        13'd2873: tone = `NM11 << 1;
        13'd2874: tone = `NM11 << 1;
        13'd2875: tone = `NM11 << 1;
        13'd2876: tone = `NM11 << 1;
        13'd2877: tone = `NM11 << 1;
        13'd2878: tone = `NM11 << 1;
        13'd2879: tone = `NM0;
        
        13'd2880: tone = `NM11 << 1;
        13'd2881: tone = `NM11 << 1;
        13'd2882: tone = `NM11 << 1;
        13'd2883: tone = `NM11 << 1;
        13'd2884: tone = `NM11 << 1;
        13'd2885: tone = `NM11 << 1;
        13'd2886: tone = `NM11 << 1;
        13'd2887: tone = `NM11 << 1;
        13'd2888: tone = `NM10 << 1;
        13'd2889: tone = `NM10 << 1;
        13'd2890: tone = `NM10 << 1;
        13'd2891: tone = `NM10 << 1;
        13'd2892: tone = `NM10 << 1;
        13'd2893: tone = `NM10 << 1;
        13'd2894: tone = `NM10 << 1;
        13'd2895: tone = `NM10 << 1;
        
        13'd2896: tone = `NM8 << 1;
        13'd2897: tone = `NM8 << 1;
        13'd2898: tone = `NM8 << 1;
        13'd2899: tone = `NM8 << 1;
        13'd2900: tone = `NM8 << 1;
        13'd2901: tone = `NM8 << 1;
        13'd2902: tone = `NM8 << 1;
        13'd2903: tone = `NM0;
        13'd2904: tone = `NM8 << 1;
        13'd2905: tone = `NM8 << 1;
        13'd2906: tone = `NM8 << 1;
        13'd2907: tone = `NM8 << 1;
        13'd2908: tone = `NM8 << 1;
        13'd2909: tone = `NM8 << 1;
        13'd2910: tone = `NM8 << 1;
        13'd2911: tone = `NM8 << 1;
        
        13'd2912: tone = `NM0;
        13'd2913: tone = `NM0;
        13'd2914: tone = `NM0;
        13'd2915: tone = `NM0;
        13'd2916: tone = `NM0;
        13'd2917: tone = `NM0;
        13'd2918: tone = `NM0;
        13'd2919: tone = `NM0;
        13'd2920: tone = `NM11 << 1;
        13'd2921: tone = `NM11 << 1;
        13'd2922: tone = `NM11 << 1;
        13'd2923: tone = `NM11 << 1;
        13'd2924: tone = `NM11 << 1;
        13'd2925: tone = `NM11 << 1;
        13'd2926: tone = `NM11 << 1;
        13'd2927: tone = `NM0;
        
        13'd2928: tone = `NM11 << 1;
        13'd2929: tone = `NM11 << 1;
        13'd2930: tone = `NM11 << 1;
        13'd2931: tone = `NM11 << 1;
        13'd2932: tone = `NM11 << 1;
        13'd2933: tone = `NM11 << 1;
        13'd2934: tone = `NM11 << 1;
        13'd2935: tone = `NM11 << 1;
        13'd2936: tone = `NM8 << 1;
        13'd2937: tone = `NM8 << 1;
        13'd2938: tone = `NM8 << 1;
        13'd2939: tone = `NM8 << 1;
        13'd2940: tone = `NM8 << 1;
        13'd2941: tone = `NM8 << 1;
        13'd2942: tone = `NM8 << 1;
        13'd2943: tone = `NM8 << 1;
        
        13'd2944: tone = `NM11 << 1;
        13'd2945: tone = `NM11 << 1;
        13'd2946: tone = `NM11 << 1;
        13'd2947: tone = `NM11 << 1;
        13'd2948: tone = `NM11 << 1;
        13'd2949: tone = `NM11 << 1;
        13'd2950: tone = `NM11 << 1;
        13'd2951: tone = `NM11 << 1;
        13'd2952: tone = `NM8 << 1;
        13'd2953: tone = `NM8 << 1;
        13'd2954: tone = `NM8 << 1;
        13'd2955: tone = `NM8 << 1;
        13'd2956: tone = `NM8 << 1;
        13'd2957: tone = `NM8 << 1;
        13'd2958: tone = `NM8 << 1;
        13'd2959: tone = `NM8 << 1;
        
        13'd2960: tone = `NM11 << 1;
        13'd2961: tone = `NM11 << 1;
        13'd2962: tone = `NM11 << 1;
        13'd2963: tone = `NM11 << 1;
        13'd2964: tone = `NM11 << 1;
        13'd2965: tone = `NM11 << 1;
        13'd2966: tone = `NM11 << 1;
        13'd2967: tone = `NM11 << 1;
        13'd2968: tone = `NM11 << 1;
        13'd2969: tone = `NM11 << 1;
        13'd2970: tone = `NM11 << 1;
        13'd2971: tone = `NM11 << 1;
        13'd2972: tone = `NM0;
        13'd2973: tone = `NM0;
        13'd2974: tone = `NM0;
        13'd2975: tone = `NM0;
        
        13'd2976: tone = `NM11 << 1;
        13'd2977: tone = `NM11 << 1;
        13'd2978: tone = `NM11 << 1;
        13'd2979: tone = `NM11 << 1;
        13'd2980: tone = `NM11 << 1;
        13'd2981: tone = `NM11 << 1;
        13'd2982: tone = `NM11 << 1;
        13'd2983: tone = `NM11 << 1;
        13'd2984: tone = `NM11 << 1;
        13'd2985: tone = `NM11 << 1;
        13'd2986: tone = `NM11 << 1;
        13'd2987: tone = `NM11 << 1;
        13'd2988: tone = `NM11 << 1;
        13'd2989: tone = `NM11 << 1;
        13'd2990: tone = `NM11 << 1;
        13'd2991: tone = `NM0;
        
        13'd2992: tone = `NM11 << 1;
        13'd2993: tone = `NM11 << 1;
        13'd2994: tone = `NM11 << 1;
        13'd2995: tone = `NM11 << 1;
        13'd2996: tone = `NM11 << 1;
        13'd2997: tone = `NM11 << 1;
        13'd2998: tone = `NM11 << 1;
        13'd2999: tone = `NM0;
        13'd3000: tone = `NM11 << 1;
        13'd3001: tone = `NM11 << 1;
        13'd3002: tone = `NM11 << 1;
        13'd3003: tone = `NM11 << 1;
        13'd3004: tone = `NM11 << 1;
        13'd3005: tone = `NM11 << 1;
        13'd3006: tone = `NM11 << 1;
        13'd3007: tone = `NM11 << 1;
        
        13'd3008: tone = `NM1 << 2;
        13'd3009: tone = `NM1 << 2;
        13'd3010: tone = `NM1 << 2;
        13'd3011: tone = `NM1 << 2;
        13'd3012: tone = `NM1 << 2;
        13'd3013: tone = `NM1 << 2;
        13'd3014: tone = `NM1 << 2;
        13'd3015: tone = `NM1 << 2;
        13'd3016: tone = `NM11 << 1;
        13'd3017: tone = `NM11 << 1;
        13'd3018: tone = `NM11 << 1;
        13'd3019: tone = `NM11 << 1;
        13'd3020: tone = `NM11 << 1;
        13'd3021: tone = `NM11 << 1;
        13'd3022: tone = `NM11 << 1;
        13'd3023: tone = `NM11 << 1;
        
        13'd3024: tone = `NM8 << 1;
        13'd3025: tone = `NM8 << 1;
        13'd3026: tone = `NM8 << 1;
        13'd3027: tone = `NM8 << 1;
        13'd3028: tone = `NM8 << 1;
        13'd3029: tone = `NM8 << 1;
        13'd3030: tone = `NM8 << 1;
        13'd3031: tone = `NM0;
        13'd3032: tone = `NM8 << 1;
        13'd3033: tone = `NM8 << 1;
        13'd3034: tone = `NM8 << 1;
        13'd3035: tone = `NM8 << 1;
        13'd3036: tone = `NM8 << 1;
        13'd3037: tone = `NM8 << 1;
        13'd3038: tone = `NM8 << 1;
        13'd3039: tone = `NM8 << 1;
        
        13'd3040: tone = `NM0;
        13'd3041: tone = `NM0;
        13'd3042: tone = `NM0;
        13'd3043: tone = `NM0;
        13'd3044: tone = `NM0;
        13'd3045: tone = `NM0;
        13'd3046: tone = `NM0;
        13'd3047: tone = `NM0;
        13'd3048: tone = `NM11 << 1;
        13'd3049: tone = `NM11 << 1;
        13'd3050: tone = `NM11 << 1;
        13'd3051: tone = `NM11 << 1;
        13'd3052: tone = `NM11 << 1;
        13'd3053: tone = `NM11 << 1;
        13'd3054: tone = `NM11 << 1;
        13'd3055: tone = `NM0;
        
        13'd3056: tone = `NM11 << 1;
        13'd3057: tone = `NM11 << 1;
        13'd3058: tone = `NM11 << 1;
        13'd3059: tone = `NM11 << 1;
        13'd3060: tone = `NM11 << 1;
        13'd3061: tone = `NM11 << 1;
        13'd3062: tone = `NM11 << 1;
        13'd3063: tone = `NM11 << 1;
        13'd3064: tone = `NM8 << 1;
        13'd3065: tone = `NM8 << 1;
        13'd3066: tone = `NM8 << 1;
        13'd3067: tone = `NM8 << 1;
        13'd3068: tone = `NM8 << 1;
        13'd3069: tone = `NM8 << 1;
        13'd3070: tone = `NM8 << 1;
        13'd3071: tone = `NM8 << 1;
        
        13'd3072: tone = `NM11 << 1;
        13'd3073: tone = `NM11 << 1;
        13'd3074: tone = `NM11 << 1;
        13'd3075: tone = `NM11 << 1;
        13'd3076: tone = `NM11 << 1;
        13'd3077: tone = `NM11 << 1;
        13'd3078: tone = `NM11 << 1;
        13'd3079: tone = `NM11 << 1;
        13'd3080: tone = `NM8 << 1;
        13'd3081: tone = `NM8 << 1;
        13'd3082: tone = `NM8 << 1;
        13'd3083: tone = `NM8 << 1;
        13'd3084: tone = `NM8 << 1;
        13'd3085: tone = `NM8 << 1;
        13'd3086: tone = `NM8 << 1;
        13'd3087: tone = `NM8 << 1;
        
        13'd3088: tone = `NM11 << 1;
        13'd3089: tone = `NM11 << 1;
        13'd3090: tone = `NM11 << 1;
        13'd3091: tone = `NM11 << 1;
        13'd3092: tone = `NM11 << 1;
        13'd3093: tone = `NM11 << 1;
        13'd3094: tone = `NM11 << 1;
        13'd3095: tone = `NM11 << 1;
        13'd3096: tone = `NM11 << 1;
        13'd3097: tone = `NM11 << 1;
        13'd3098: tone = `NM11 << 1;
        13'd3099: tone = `NM11 << 1;
        13'd3100: tone = `NM0;
        13'd3101: tone = `NM0;
        13'd3102: tone = `NM0;
        13'd3103: tone = `NM0;
        
        13'd3104: tone = `NM11 << 1;
        13'd3105: tone = `NM11 << 1;
        13'd3106: tone = `NM11 << 1;
        13'd3107: tone = `NM11 << 1;
        13'd3108: tone = `NM11 << 1;
        13'd3109: tone = `NM11 << 1;
        13'd3110: tone = `NM11 << 1;
        13'd3111: tone = `NM11 << 1;
        13'd3112: tone = `NM11 << 1;
        13'd3113: tone = `NM11 << 1;
        13'd3114: tone = `NM11 << 1;
        13'd3115: tone = `NM11 << 1;
        13'd3116: tone = `NM11 << 1;
        13'd3117: tone = `NM11 << 1;
        13'd3118: tone = `NM11 << 1;
        13'd3119: tone = `NM0;
        
        13'd3120: tone = `NM11 << 1;
        13'd3121: tone = `NM11 << 1;
        13'd3122: tone = `NM11 << 1;
        13'd3123: tone = `NM11 << 1;
        13'd3124: tone = `NM11 << 1;
        13'd3125: tone = `NM11 << 1;
        13'd3126: tone = `NM11 << 1;
        13'd3127: tone = `NM0;
        13'd3128: tone = `NM11 << 1;
        13'd3129: tone = `NM11 << 1;
        13'd3130: tone = `NM11 << 1;
        13'd3131: tone = `NM11 << 1;
        13'd3132: tone = `NM11 << 1;
        13'd3133: tone = `NM11 << 1;
        13'd3134: tone = `NM11 << 1;
        13'd3135: tone = `NM0;
        
        13'd3136: tone = `NM11 << 1;
        13'd3137: tone = `NM11 << 1;
        13'd3138: tone = `NM11 << 1;
        13'd3139: tone = `NM11 << 1;
        13'd3140: tone = `NM11 << 1;
        13'd3141: tone = `NM11 << 1;
        13'd3142: tone = `NM11 << 1;
        13'd3143: tone = `NM0;
        13'd3144: tone = `NM10 << 1;
        13'd3145: tone = `NM10 << 1;
        13'd3146: tone = `NM10 << 1;
        13'd3147: tone = `NM10 << 1;
        13'd3148: tone = `NM10 << 1;
        13'd3149: tone = `NM10 << 1;
        13'd3150: tone = `NM10 << 1;
        13'd3151: tone = `NM0;
        
        13'd3152: tone = `NM8 << 1;
        13'd3153: tone = `NM8 << 1;
        13'd3154: tone = `NM8 << 1;
        13'd3155: tone = `NM8 << 1;
        13'd3156: tone = `NM8 << 1;
        13'd3157: tone = `NM8 << 1;
        13'd3158: tone = `NM8 << 1;
        13'd3159: tone = `NM0;
        13'd3160: tone = `NM8 << 1;
        13'd3161: tone = `NM8 << 1;
        13'd3162: tone = `NM8 << 1;
        13'd3163: tone = `NM8 << 1;
        13'd3164: tone = `NM8 << 1;
        13'd3165: tone = `NM8 << 1;
        13'd3166: tone = `NM8 << 1;
        13'd3167: tone = `NM8 << 1;
        
        13'd3168: tone = `NM0;
        13'd3169: tone = `NM0;
        13'd3170: tone = `NM0;
        13'd3171: tone = `NM0;
        13'd3172: tone = `NM0;
        13'd3173: tone = `NM0;
        13'd3174: tone = `NM0;
        13'd3175: tone = `NM0;
        13'd3176: tone = `NM6 << 1;
        13'd3177: tone = `NM6 << 1;
        13'd3178: tone = `NM6 << 1;
        13'd3179: tone = `NM6 << 1;
        13'd3180: tone = `NM6 << 1;
        13'd3181: tone = `NM6 << 1;
        13'd3182: tone = `NM6 << 1;
        13'd3183: tone = `NM0;
        
        13'd3184: tone = `NM6 << 1;
        13'd3185: tone = `NM6 << 1;
        13'd3186: tone = `NM6 << 1;
        13'd3187: tone = `NM6 << 1;
        13'd3188: tone = `NM6 << 1;
        13'd3189: tone = `NM6 << 1;
        13'd3190: tone = `NM6 << 1;
        13'd3191: tone = `NM6 << 1;
        13'd3192: tone = `NM8 << 1;
        13'd3193: tone = `NM8 << 1;
        13'd3194: tone = `NM8 << 1;
        13'd3195: tone = `NM8 << 1;
        13'd3196: tone = `NM8 << 1;
        13'd3197: tone = `NM8 << 1;
        13'd3198: tone = `NM8 << 1;
        13'd3199: tone = `NM8 << 1;
        
        13'd3200: tone = `NM0;
        13'd3201: tone = `NM0;
        13'd3202: tone = `NM0;
        13'd3203: tone = `NM0;
        13'd3204: tone = `NM0;
        13'd3205: tone = `NM0;
        13'd3206: tone = `NM0;
        13'd3207: tone = `NM0;
        13'd3208: tone = `NM6 << 1;
        13'd3209: tone = `NM6 << 1;
        13'd3210: tone = `NM6 << 1;
        13'd3211: tone = `NM6 << 1;
        13'd3212: tone = `NM6 << 1;
        13'd3213: tone = `NM6 << 1;
        13'd3214: tone = `NM6 << 1;
        13'd3215: tone = `NM0;
        
        13'd3216: tone = `NM6 << 1;
        13'd3217: tone = `NM6 << 1;
        13'd3218: tone = `NM6 << 1;
        13'd3219: tone = `NM6 << 1;
        13'd3220: tone = `NM6 << 1;
        13'd3221: tone = `NM6 << 1;
        13'd3222: tone = `NM6 << 1;
        13'd3223: tone = `NM0;
        13'd3224: tone = `NM8 << 1;
        13'd3225: tone = `NM8 << 1;
        13'd3226: tone = `NM8 << 1;
        13'd3227: tone = `NM8 << 1;
        13'd3228: tone = `NM8 << 1;
        13'd3229: tone = `NM8 << 1;
        13'd3230: tone = `NM8 << 1;
        13'd3231: tone = `NM8 << 1;
        
        13'd3232: tone = `NM0;
        13'd3233: tone = `NM0;
        13'd3234: tone = `NM0;
        13'd3235: tone = `NM0;
        13'd3236: tone = `NM0;
        13'd3237: tone = `NM0;
        13'd3238: tone = `NM0;
        13'd3239: tone = `NM0;
        13'd3240: tone = `NM8 << 1;
        13'd3241: tone = `NM8 << 1;
        13'd3242: tone = `NM8 << 1;
        13'd3243: tone = `NM8 << 1;
        13'd3244: tone = `NM8 << 1;
        13'd3245: tone = `NM8 << 1;
        13'd3246: tone = `NM8 << 1;
        13'd3247: tone = `NM0;
        
        13'd3248: tone = `NM8 << 1;
        13'd3249: tone = `NM8 << 1;
        13'd3250: tone = `NM8 << 1;
        13'd3251: tone = `NM8 << 1;
        13'd3252: tone = `NM8 << 1;
        13'd3253: tone = `NM8 << 1;
        13'd3254: tone = `NM8 << 1;
        13'd3255: tone = `NM8 << 1;
        13'd3256: tone = `NM11 << 1;
        13'd3257: tone = `NM11 << 1;
        13'd3258: tone = `NM11 << 1;
        13'd3259: tone = `NM11 << 1;
        13'd3260: tone = `NM11 << 1;
        13'd3261: tone = `NM11 << 1;
        13'd3262: tone = `NM11 << 1;
        13'd3263: tone = `NM11 << 1;
        
        13'd3264: tone = `NM0;
        13'd3265: tone = `NM0;
        13'd3266: tone = `NM0;
        13'd3267: tone = `NM0;
        13'd3268: tone = `NM0;
        13'd3269: tone = `NM0;
        13'd3270: tone = `NM0;
        13'd3271: tone = `NM0;
        13'd3272: tone = `NM8 << 1;
        13'd3273: tone = `NM8 << 1;
        13'd3274: tone = `NM8 << 1;
        13'd3275: tone = `NM8 << 1;
        13'd3276: tone = `NM8 << 1;
        13'd3277: tone = `NM8 << 1;
        13'd3278: tone = `NM8 << 1;
        13'd3279: tone = `NM0;
        
        13'd3280: tone = `NM8 << 1;
        13'd3281: tone = `NM8 << 1;
        13'd3282: tone = `NM8 << 1;
        13'd3283: tone = `NM8 << 1;
        13'd3284: tone = `NM8 << 1;
        13'd3285: tone = `NM8 << 1;
        13'd3286: tone = `NM8 << 1;
        13'd3287: tone = `NM8 << 1;
        13'd3288: tone = `NM11 << 1;
        13'd3289: tone = `NM11 << 1;
        13'd3290: tone = `NM11 << 1;
        13'd3291: tone = `NM11 << 1;
        13'd3292: tone = `NM11 << 1;
        13'd3293: tone = `NM11 << 1;
        13'd3294: tone = `NM11 << 1;
        13'd3295: tone = `NM11 << 1;
        
        13'd3296: tone = `NM11 << 1;
        13'd3297: tone = `NM11 << 1;
        13'd3298: tone = `NM11 << 1;
        13'd3299: tone = `NM11 << 1;
        13'd3300: tone = `NM11 << 1;
        13'd3301: tone = `NM11 << 1;
        13'd3302: tone = `NM11 << 1;
        13'd3303: tone = `NM0;
        13'd3304: tone = `NM11 << 1;
        13'd3305: tone = `NM11 << 1;
        13'd3306: tone = `NM11 << 1;
        13'd3307: tone = `NM11 << 1;
        13'd3308: tone = `NM11 << 1;
        13'd3309: tone = `NM11 << 1;
        13'd3310: tone = `NM11 << 1;
        13'd3311: tone = `NM11 << 1;
        
        13'd3312: tone = `NM1 << 2;
        13'd3313: tone = `NM1 << 2;
        13'd3314: tone = `NM1 << 2;
        13'd3315: tone = `NM1 << 2;
        13'd3316: tone = `NM1 << 2;
        13'd3317: tone = `NM1 << 2;
        13'd3318: tone = `NM1 << 2;
        13'd3319: tone = `NM1 << 2;
        13'd3320: tone = `NM11 << 1;
        13'd3321: tone = `NM11 << 1;
        13'd3322: tone = `NM11 << 1;
        13'd3323: tone = `NM11 << 1;
        13'd3324: tone = `NM11 << 1;
        13'd3325: tone = `NM11 << 1;
        13'd3326: tone = `NM11 << 1;
        13'd3327: tone = `NM11 << 1;
        
        13'd3328: tone = `NM11 << 1;
        13'd3329: tone = `NM11 << 1;
        13'd3330: tone = `NM11 << 1;
        13'd3331: tone = `NM11 << 1;
        13'd3332: tone = `NM11 << 1;
        13'd3333: tone = `NM11 << 1;
        13'd3334: tone = `NM11 << 1;
        13'd3335: tone = `NM11 << 1;
        13'd3336: tone = `NM11 << 1;
        13'd3337: tone = `NM11 << 1;
        13'd3338: tone = `NM11 << 1;
        13'd3339: tone = `NM11 << 1;
        13'd3340: tone = `NM11 << 1;
        13'd3341: tone = `NM11 << 1;
        13'd3342: tone = `NM11 << 1;
        13'd3343: tone = `NM11 << 1;
        // 000
     
        13'd3344: tone = `NM0;
        13'd3345: tone = `NM0;
        13'd3346: tone = `NM0;
        13'd3347: tone = `NM0;
        13'd3348: tone = `NM0;
        13'd3349: tone = `NM0;
        13'd3350: tone = `NM0;
        13'd3351: tone = `NM0;
        13'd3352: tone = `NM0;
        13'd3353: tone = `NM0;
        13'd3354: tone = `NM0;
        13'd3355: tone = `NM0;
        13'd3356: tone = `NM0;
        13'd3357: tone = `NM0;
        13'd3358: tone = `NM0;
        13'd3359: tone = `NM0;
        
       13'd3360: tone = `NM8 << 1;
        13'd3361: tone = `NM8 << 1;
        13'd3362: tone = `NM8 << 1;
        13'd3363: tone = `NM8 << 1;
        13'd3364: tone = `NM8 << 1;
        13'd3365: tone = `NM8 << 1;
        13'd3366: tone = `NM8 << 1;
        13'd3367: tone = `NM8 << 1;
        13'd3368: tone = `NM8 << 1;
        13'd3369: tone = `NM8 << 1;
        13'd3370: tone = `NM8 << 1;
        13'd3371: tone = `NM8 << 1;
        13'd3372: tone = `NM8 << 1;
        13'd3373: tone = `NM8 << 1;
        13'd3374: tone = `NM8 << 1;
        13'd3375: tone = `NM8 << 1;
        
        13'd3376: tone = `NM8 << 1;
        13'd3377: tone = `NM8 << 1;
        13'd3378: tone = `NM8 << 1;
        13'd3379: tone = `NM8 << 1;
        13'd3380: tone = `NM8 << 1;
        13'd3381: tone = `NM8 << 1;
        13'd3382: tone = `NM8 << 1;
        13'd3383: tone = `NM8 << 1;
        13'd3384: tone = `NM8 << 1;
        13'd3385: tone = `NM8 << 1;
        13'd3386: tone = `NM8 << 1;
        13'd3387: tone = `NM8 << 1;
        13'd3388: tone = `NM8 << 1;
        13'd3389: tone = `NM8 << 1;
        13'd3390: tone = `NM8 << 1;
        13'd3391: tone = `NM0;
        
        13'd3392: tone = `NM8 << 1;
        13'd3393: tone = `NM8 << 1;
        13'd3394: tone = `NM8 << 1;
        13'd3395: tone = `NM8 << 1;
        13'd3396: tone = `NM8 << 1;
        13'd3397: tone = `NM8 << 1;
        13'd3398: tone = `NM8 << 1;
        13'd3399: tone = `NM8 << 1;
        13'd3400: tone = `NM8 << 1;
        13'd3401: tone = `NM8 << 1;
        13'd3402: tone = `NM8 << 1;
        13'd3403: tone = `NM8 << 1;
        13'd3404: tone = `NM8 << 1;
        13'd3405: tone = `NM8 << 1;
        13'd3406: tone = `NM8 << 1;
        13'd3407: tone = `NM8 << 1;
        
        13'd3408: tone = `NM8 << 1;
        13'd3409: tone = `NM8 << 1;
        13'd3410: tone = `NM8 << 1;
        13'd3411: tone = `NM8 << 1;
        13'd3412: tone = `NM8 << 1;
        13'd3413: tone = `NM8 << 1;
        13'd3414: tone = `NM8 << 1;
        13'd3415: tone = `NM8 << 1;
        13'd3416: tone = `NM8 << 1;
        13'd3417: tone = `NM8 << 1;
        13'd3418: tone = `NM8 << 1;
        13'd3419: tone = `NM8 << 1;
        13'd3420: tone = `NM8 << 1;
        13'd3421: tone = `NM8 << 1;
        13'd3422: tone = `NM8 << 1;
        13'd3423: tone = `NM0;
        
        13'd3424: tone = `NM8 << 1;
        13'd3425: tone = `NM8 << 1;
        13'd3426: tone = `NM8 << 1;
        13'd3427: tone = `NM8 << 1;
        13'd3428: tone = `NM8 << 1;
        13'd3429: tone = `NM8 << 1;
        13'd3430: tone = `NM8 << 1;
        13'd3431: tone = `NM8 << 1;
        13'd3432: tone = `NM8 << 1;
        13'd3433: tone = `NM8 << 1;
        13'd3434: tone = `NM8 << 1;
        13'd3435: tone = `NM8 << 1;
        13'd3436: tone = `NM8 << 1;
        13'd3437: tone = `NM8 << 1;
        13'd3438: tone = `NM8 << 1;
        13'd3439: tone = `NM8 << 1;
        
        13'd3440: tone = `NM8 << 1;
        13'd3441: tone = `NM8 << 1;
        13'd3442: tone = `NM8 << 1;
        13'd3443: tone = `NM8 << 1;
        13'd3444: tone = `NM8 << 1;
        13'd3445: tone = `NM8 << 1;
        13'd3446: tone = `NM8 << 1;
        13'd3447: tone = `NM8 << 1;
        13'd3448: tone = `NM8 << 1;
        13'd3449: tone = `NM8 << 1;
        13'd3450: tone = `NM8 << 1;
        13'd3451: tone = `NM8 << 1;
        13'd3452: tone = `NM8 << 1;
        13'd3453: tone = `NM8 << 1;
        13'd3454: tone = `NM8 << 1;
        13'd3455: tone = `NM8 << 1;

        13'd3456: tone = `NM0;
        13'd3457: tone = `NM0;
        13'd3458: tone = `NM0;
        13'd3459: tone = `NM0;
        13'd3460: tone = `NM0;
        13'd3461: tone = `NM0;
        13'd3462: tone = `NM0;
        13'd3463: tone = `NM0;
		default : tone = `NM0;
    
        

	endcase
end

endmodule